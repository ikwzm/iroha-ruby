// Generated from iroha-0.1.0.

module fadd(clk, rst_n, i_valid, z_out, a_in, b_in, sub);
  input clk;
  input rst_n;
  input i_valid;
  output [31:0] z_out;
  input [31:0] a_in;
  input [31:0] b_in;
  input sub;
  reg [31:0] z_out;

  // State decls
  reg st_1_1;
  reg st_1_2;
  reg st_1_3;
  reg st_1_4;
  reg st_1_5;
  reg st_1_6;
  reg st_1_7;
  reg st_1_8;
  // State vars
  // Registers
  wire  [0:0] start;
  reg  [22:0] stage1_a_fraction;
  reg  [7:0] stage1_a_exponent;
  reg  stage1_a_sign;
  reg  [22:0] stage1_b_fraction;
  reg  [7:0] stage1_b_exponent;
  reg  stage1_b_sign;
  reg  stage1_sub;
  reg  stage2_sub;
  reg  stage2_b_gt_a;
  reg  [23:0] stage2_l_fraction;
  reg  [7:0] stage2_l_exponent;
  reg  stage2_l_sign;
  reg  [23:0] stage2_s_fraction;
  reg  [7:0] stage2_s_exponent;
  reg  stage2_s_sign;
  reg  stage2_a_is_zero;
  reg  stage2_a_is_inf;
  reg  stage2_a_is_nan;
  reg  stage2_b_is_zero;
  reg  stage2_b_is_inf;
  reg  stage2_b_is_nan;
  reg  stage3_sub;
  reg  stage3_b_gt_a;
  reg  stage3_op_sub;
  reg  [7:0] stage3_diff_exponent;
  reg  [0:0] stage3_t_sign;
  reg  [7:0] stage3_t_exponent;
  reg  [23:0] stage3_l_fraction;
  reg  [23:0] stage3_s_fraction;
  reg  stage3_a_is_zero;
  reg  stage3_a_is_inf;
  reg  stage3_a_is_nan;
  reg  stage3_b_is_zero;
  reg  stage3_b_is_inf;
  reg  stage3_b_is_nan;
  reg  stage4_sub;
  reg  stage4_b_gt_a;
  reg  stage4_op_sub;
  reg  [0:0] stage4_t_sign;
  reg  [7:0] stage4_t_exponent;
  reg  [27:0] stage4_l_fraction;
  reg  [27:0] stage4_s_fraction;
  reg  stage4_a_is_zero;
  reg  stage4_a_is_inf;
  reg  stage4_a_is_nan;
  reg  stage4_b_is_zero;
  reg  stage4_b_is_inf;
  reg  stage4_b_is_nan;
  reg  stage5_sub;
  reg  stage5_b_gt_a;
  reg  [0:0] stage5_t_sign;
  reg  [7:0] stage5_t_exponent;
  reg  [27:0] stage5_t_fraction;
  reg  stage5_a_is_zero;
  reg  stage5_a_is_inf;
  reg  stage5_a_is_nan;
  reg  stage5_b_is_zero;
  reg  stage5_b_is_inf;
  reg  stage5_b_is_nan;
  reg  stage6_sub;
  reg  stage6_b_gt_a;
  reg  [0:0] stage6_t_sign;
  reg  signed [8:0] stage6_t_exponent;
  reg  [27:0] stage6_t_fraction;
  reg  stage6_a_is_zero;
  reg  stage6_a_is_inf;
  reg  stage6_a_is_nan;
  reg  stage6_b_is_zero;
  reg  stage6_b_is_inf;
  reg  stage6_b_is_nan;
  reg  stage7_sub;
  reg  stage7_b_gt_a;
  reg  [0:0] stage7_t_sign;
  reg  signed [8:0] stage7_t_exponent;
  reg  [23:0] stage7_t_fraction;
  reg  stage7_a_is_zero;
  reg  stage7_a_is_inf;
  reg  stage7_a_is_nan;
  reg  stage7_b_is_zero;
  reg  stage7_b_is_inf;
  reg  stage7_b_is_nan;
  wire  [31:0] stage1_a_data_in;
  wire  [22:0] stage1_a_fraction_in;
  wire  [7:0] stage1_a_exponent_in;
  wire  [31:0] stage1_b_data_in;
  wire  [22:0] stage1_b_fraction_in;
  wire  [7:0] stage1_b_exponent_in;
  wire  stage2_a_exponent_is_all_1;
  wire  stage2_a_exponent_is_all_0;
  wire  stage2_a_fraction_is_all_0;
  wire  stage2_a_fraction_is_not_0;
  wire  [0:0] stage2_a_fraction_msb;
  wire  [23:0] stage2_a_fraction_in;
  wire  [7:0] stage2_a_exponent_in;
  wire  [0:0] stage2_a_sign_in;
  wire  stage2_b_exponent_is_all_1;
  wire  stage2_b_exponent_is_all_0;
  wire  stage2_b_fraction_is_all_0;
  wire  stage2_b_fraction_is_not_0;
  wire  [0:0] stage2_b_fraction_msb;
  wire  [23:0] stage2_b_fraction_in;
  wire  [7:0] stage2_b_exponent_in;
  wire  [0:0] stage2_b_sign_in;
  wire  [30:0] stage2_a_abs_data;
  wire  [30:0] stage2_b_abs_data;
  wire  stage2_b_gt_a_125;
  wire  stage3_sub_xor_l_sign;
  wire  [51:0] stage4_shift_fractions_0;
  wire  [51:0] stage4_shift_fractions_1;
  wire  [51:0] stage4_shift_fractions_2;
  wire  [51:0] stage4_shift_fractions_3;
  wire  [51:0] stage4_shift_fractions_4;
  wire  [51:0] stage4_shift_fractions_5;
  wire  [0:0] anon_141;
  wire  [50:0] anon_142;
  wire  [51:0] anon_143;
  wire  [0:0] anon_149;
  wire  [49:0] anon_150;
  wire  [51:0] anon_151;
  wire  [0:0] anon_157;
  wire  [47:0] anon_158;
  wire  [51:0] anon_159;
  wire  [0:0] anon_165;
  wire  [43:0] anon_166;
  wire  [51:0] anon_167;
  wire  [0:0] anon_173;
  wire  [35:0] anon_174;
  wire  [51:0] anon_175;
  wire  [26:0] stage4_s_fraction_data;
  wire  [27:0] stage4_s_fraction_181;
  wire  [24:0] stage4_s_sticky_data;
  wire  [0:0] stage4_s_sticky;
  wire  stage4_s_under;
  wire  anon_191;
  wire  [27:0] stage5_add_s_fraction;
  wire  [27:0] stage5_sub_s_fraction;
  wire  [27:0] stage5_s_fraction;
  wire  [27:0] anon_196;
  wire  [4:0] stage6_shift;
  wire  [0:0] stage6_shift_flag_0;
  wire  [0:0] stage6_shift_flag_1;
  wire  [0:0] stage6_shift_flag_2;
  wire  [0:0] stage6_shift_flag_3;
  wire  [0:0] stage6_shift_flag_4;
  wire  [27:0] stage6_fraction_data_0;
  wire  [27:0] stage6_fraction_data_1;
  wire  [27:0] stage6_fraction_data_2;
  wire  [27:0] stage6_fraction_data_3;
  wire  [27:0] stage6_fraction_data_4;
  wire  [27:0] stage6_fraction_data_5;
  wire  signed [8:0] stage6_exponent_data;
  wire  [15:0] anon_214;
  wire  [11:0] anon_218;
  wire  [27:0] anon_219;
  wire  [7:0] anon_223;
  wire  [19:0] anon_227;
  wire  [27:0] anon_228;
  wire  [3:0] anon_232;
  wire  [23:0] anon_236;
  wire  [27:0] anon_237;
  wire  [1:0] anon_241;
  wire  [25:0] anon_245;
  wire  [27:0] anon_246;
  wire  [0:0] anon_250;
  wire  [26:0] anon_254;
  wire  [27:0] anon_255;
  wire  signed [8:0] anon_257;
  wire  [23:0] stage7_fraction_data;
  wire  [0:0] stage7_ulp;
  wire  [0:0] stage7_uulp1;
  wire  [0:0] stage7_uulp2;
  wire  [0:0] stage7_uulp3;
  wire  [0:0] stage7_uulp4;
  wire  [0:0] stage7_increment;
  wire  [0:0] anon_278;
  wire  [0:0] anon_279;
  wire  [0:0] anon_280;
  wire  anon_281;
  wire  [0:0] anon_282;
  wire  stage8_set_nan;
  wire  stage8_set_inf;
  wire  stage8_set_zero;
  wire  anon_293;
  wire  anon_294;
  wire  anon_295;
  wire  anon_296;
  wire  anon_297;
  wire  [0:0] stage8_fraction_msb;
  wire  [22:0] stage8_fraction_in;
  wire  [7:0] stage8_exponent_in;
  wire  [0:0] stage8_sign_in;
  wire  stage8_exp_natural;
  wire  stage8_exp_underflow;
  wire  stage8_exp_overflow;
  wire  anon_312;
  wire  [0:0] anon_313;
  wire  anon_315;
  wire  [22:0] stage8_fraction_i1;
  wire  [7:0] stage8_exponent_i1;
  wire  [0:0] stage8_sign_i1;
  wire  [22:0] stage8_fraction_i2;
  wire  [7:0] stage8_exponent_i2;
  wire  [0:0] stage8_sign_i2;
  wire  [22:0] stage8_fraction_i3;
  wire  [7:0] stage8_exponent_i3;
  wire  [0:0] stage8_sign_i3;
  wire  [22:0] stage8_fraction_i4;
  wire  [7:0] stage8_exponent_i4;
  wire  [0:0] stage8_sign_i4;
  wire  [22:0] stage8_fraction_o;
  wire  [7:0] stage8_exponent_o;
  wire  [0:0] stage8_sign_o;
  wire  [31:0] stage8_result;
  // Resources
  // eq:18
  wire [7:0] eq_18_s0;
  assign eq_18_s0 = stage1_a_exponent;
  wire [7:0] eq_18_s1;
  assign eq_18_s1 = 8'd255;
  wire eq_18_d0;
  assign eq_18_d0 = eq_18_s0 == eq_18_s1;
  // eq:19
  wire [7:0] eq_19_s0;
  assign eq_19_s0 = stage1_a_exponent;
  wire [7:0] eq_19_s1;
  assign eq_19_s1 = 8'd0;
  wire eq_19_d0;
  assign eq_19_d0 = eq_19_s0 == eq_19_s1;
  // eq:20
  wire [22:0] eq_20_s0;
  assign eq_20_s0 = stage1_a_fraction;
  wire [22:0] eq_20_s1;
  assign eq_20_s1 = 23'd0;
  wire eq_20_d0;
  assign eq_20_d0 = eq_20_s0 == eq_20_s1;
  // eq:29
  wire [7:0] eq_29_s0;
  assign eq_29_s0 = stage1_b_exponent;
  wire [7:0] eq_29_s1;
  assign eq_29_s1 = 8'd255;
  wire eq_29_d0;
  assign eq_29_d0 = eq_29_s0 == eq_29_s1;
  // eq:30
  wire [7:0] eq_30_s0;
  assign eq_30_s0 = stage1_b_exponent;
  wire [7:0] eq_30_s1;
  assign eq_30_s1 = 8'd0;
  wire eq_30_d0;
  assign eq_30_d0 = eq_30_s0 == eq_30_s1;
  // eq:31
  wire [22:0] eq_31_s0;
  assign eq_31_s0 = stage1_b_fraction;
  wire [22:0] eq_31_s1;
  assign eq_31_s1 = 23'd0;
  wire eq_31_d0;
  assign eq_31_d0 = eq_31_s0 == eq_31_s1;
  // gt:42
  wire [30:0] gt_42_s0;
  assign gt_42_s0 = stage2_b_abs_data;
  wire [30:0] gt_42_s1;
  assign gt_42_s1 = stage2_a_abs_data;
  wire gt_42_d0;
  assign gt_42_d0 = gt_42_s0 > gt_42_s1;
  // sub:54
  wire [7:0] sub_54_s0;
  assign sub_54_s0 = stage2_l_exponent;
  wire [7:0] sub_54_s1;
  assign sub_54_s1 = stage2_s_exponent;
  wire [7:0] sub_54_d0;
  assign sub_54_d0 = sub_54_s0 - sub_54_s1;
  // gte:87
  wire [7:0] gte_87_s0;
  assign gte_87_s0 = stage3_diff_exponent;
  wire [5:0] gte_87_s1;
  assign gte_87_s1 = 6'd28;
  wire gte_87_d0;
  assign gte_87_d0 = gte_87_s0 >= gte_87_s1;
  // eq:90
  wire [24:0] eq_90_s0;
  assign eq_90_s0 = stage4_s_sticky_data;
  wire [24:0] eq_90_s1;
  assign eq_90_s1 = 25'd0;
  wire eq_90_d0;
  assign eq_90_d0 = eq_90_s0 == eq_90_s1;
  // add:108
  wire [27:0] add_108_s0;
  assign add_108_s0 = anon_196;
  wire [27:0] add_108_s1;
  assign add_108_s1 = 28'd1;
  wire [27:0] add_108_d0;
  assign add_108_d0 = add_108_s0 + add_108_s1;
  // add:110
  wire [27:0] add_110_s0;
  assign add_110_s0 = stage4_l_fraction;
  wire [27:0] add_110_s1;
  assign add_110_s1 = stage5_s_fraction;
  wire [27:0] add_110_d0;
  assign add_110_d0 = add_110_s0 + add_110_s1;
  // eq:123
  wire [15:0] eq_123_s0;
  assign eq_123_s0 = anon_214;
  wire [15:0] eq_123_s1;
  assign eq_123_s1 = 16'd0;
  wire [0:0] eq_123_d0;
  assign eq_123_d0 = eq_123_s0 == eq_123_s1;
  // eq:128
  wire [7:0] eq_128_s0;
  assign eq_128_s0 = anon_223;
  wire [7:0] eq_128_s1;
  assign eq_128_s1 = 8'd0;
  wire [0:0] eq_128_d0;
  assign eq_128_d0 = eq_128_s0 == eq_128_s1;
  // eq:133
  wire [3:0] eq_133_s0;
  assign eq_133_s0 = anon_232;
  wire [3:0] eq_133_s1;
  assign eq_133_s1 = 4'd0;
  wire [0:0] eq_133_d0;
  assign eq_133_d0 = eq_133_s0 == eq_133_s1;
  // eq:138
  wire [1:0] eq_138_s0;
  assign eq_138_s0 = anon_241;
  wire [1:0] eq_138_s1;
  assign eq_138_s1 = 2'd0;
  wire [0:0] eq_138_d0;
  assign eq_138_d0 = eq_138_s0 == eq_138_s1;
  // eq:143
  wire [0:0] eq_143_s0;
  assign eq_143_s0 = anon_250;
  wire [0:0] eq_143_s1;
  assign eq_143_s1 = 1'd0;
  wire [0:0] eq_143_d0;
  assign eq_143_d0 = eq_143_s0 == eq_143_s1;
  // sub:148
  wire [7:0] sub_148_s0;
  assign sub_148_s0 = stage5_t_exponent;
  wire [4:0] sub_148_s1;
  assign sub_148_s1 = stage6_shift;
  wire signed [8:0] sub_148_d0;
  assign sub_148_d0 = sub_148_s0 - sub_148_s1;
  // add:149
  wire signed [8:0] add_149_s0;
  assign add_149_s0 = anon_257;
  wire [0:0] add_149_s1;
  assign add_149_s1 = 1'd1;
  wire signed [8:0] add_149_d0;
  assign add_149_d0 = add_149_s0 + add_149_s1;
  // add:170
  wire [23:0] add_170_s0;
  assign add_170_s0 = stage7_fraction_data;
  wire [0:0] add_170_s1;
  assign add_170_s1 = stage7_increment;
  wire [23:0] add_170_d0;
  assign add_170_d0 = add_170_s0 + add_170_s1;
  // eq:171
  wire [23:0] eq_171_s0;
  assign eq_171_s0 = stage7_fraction_data;
  wire [23:0] eq_171_s1;
  assign eq_171_s1 = 24'd16777215;
  wire eq_171_d0;
  assign eq_171_d0 = eq_171_s0 == eq_171_s1;
  // add:173
  wire signed [8:0] add_173_s0;
  assign add_173_s0 = stage6_t_exponent;
  wire [0:0] add_173_s1;
  assign add_173_s1 = anon_282;
  wire signed [8:0] add_173_d0;
  assign add_173_d0 = add_173_s0 + add_173_s1;
  // gt:194
  wire signed [8:0] gt_194_s0;
  assign gt_194_s0 = stage7_t_exponent;
  wire signed [8:0] gt_194_s1;
  assign gt_194_s1 = 9'd0;
  wire gt_194_d0;
  assign gt_194_d0 = gt_194_s0 > gt_194_s1;
  // gte:198
  wire signed [8:0] gte_198_s0;
  assign gte_198_s0 = stage7_t_exponent;
  wire signed [8:0] gte_198_s1;
  assign gte_198_s1 = 9'd255;
  wire gte_198_d0;
  assign gte_198_d0 = gte_198_s0 >= gte_198_s1;
  // Insn wires
  wire  [0:0] insn_o_1_9_0;
  wire  insn_o_1_10_0;
  wire  [31:0] insn_o_1_11_0;
  wire  [22:0] insn_o_1_12_0;
  wire  [7:0] insn_o_1_13_0;
  wire  insn_o_1_14_0;
  wire  [22:0] insn_o_1_15_0;
  wire  [7:0] insn_o_1_16_0;
  wire  [31:0] insn_o_1_17_0;
  wire  [22:0] insn_o_1_18_0;
  wire  [7:0] insn_o_1_19_0;
  wire  insn_o_1_20_0;
  wire  [22:0] insn_o_1_21_0;
  wire  [7:0] insn_o_1_22_0;
  wire  insn_o_1_23_0;
  wire  insn_o_1_24_0;
  wire  insn_o_1_25_0;
  wire  insn_o_1_26_0;
  wire  [0:0] insn_o_1_27_0;
  wire  [23:0] insn_o_1_28_0;
  wire  [7:0] insn_o_1_29_0;
  wire  [0:0] insn_o_1_30_0;
  wire  insn_o_1_31_0;
  wire  insn_o_1_32_0;
  wire  insn_o_1_33_0;
  wire  insn_o_1_34_0;
  wire  insn_o_1_35_0;
  wire  insn_o_1_36_0;
  wire  insn_o_1_37_0;
  wire  [0:0] insn_o_1_38_0;
  wire  [23:0] insn_o_1_39_0;
  wire  [7:0] insn_o_1_40_0;
  wire  [0:0] insn_o_1_41_0;
  wire  insn_o_1_42_0;
  wire  insn_o_1_43_0;
  wire  insn_o_1_44_0;
  wire  [30:0] insn_o_1_45_0;
  wire  [30:0] insn_o_1_46_0;
  wire  insn_o_1_47_0;
  wire  [23:0] insn_o_1_48_0;
  wire  [7:0] insn_o_1_49_0;
  wire  insn_o_1_50_0;
  wire  [23:0] insn_o_1_51_0;
  wire  [7:0] insn_o_1_52_0;
  wire  insn_o_1_53_0;
  wire  insn_o_1_54_0;
  wire  insn_o_1_55_0;
  wire  insn_o_1_56_0;
  wire  [0:0] insn_o_1_57_0;
  wire  insn_o_1_58_0;
  wire  [7:0] insn_o_1_59_0;
  wire  [7:0] insn_o_1_60_0;
  wire  [23:0] insn_o_1_61_0;
  wire  [23:0] insn_o_1_62_0;
  wire  insn_o_1_63_0;
  wire  insn_o_1_64_0;
  wire  insn_o_1_65_0;
  wire  insn_o_1_66_0;
  wire  insn_o_1_67_0;
  wire  insn_o_1_68_0;
  wire  insn_o_1_69_0;
  wire  insn_o_1_70_0;
  wire  [51:0] insn_o_1_71_0;
  wire  [0:0] insn_o_1_72_0;
  wire  [50:0] insn_o_1_73_0;
  wire  [51:0] insn_o_1_74_0;
  wire  [51:0] insn_o_1_75_0;
  wire  [0:0] insn_o_1_76_0;
  wire  [49:0] insn_o_1_77_0;
  wire  [51:0] insn_o_1_78_0;
  wire  [51:0] insn_o_1_79_0;
  wire  [0:0] insn_o_1_80_0;
  wire  [47:0] insn_o_1_81_0;
  wire  [51:0] insn_o_1_82_0;
  wire  [51:0] insn_o_1_83_0;
  wire  [0:0] insn_o_1_84_0;
  wire  [43:0] insn_o_1_85_0;
  wire  [51:0] insn_o_1_86_0;
  wire  [51:0] insn_o_1_87_0;
  wire  [0:0] insn_o_1_88_0;
  wire  [35:0] insn_o_1_89_0;
  wire  [51:0] insn_o_1_90_0;
  wire  [51:0] insn_o_1_91_0;
  wire  insn_o_1_92_0;
  wire  [26:0] insn_o_1_93_0;
  wire  [24:0] insn_o_1_94_0;
  wire  insn_o_1_95_0;
  wire  [0:0] insn_o_1_96_0;
  wire  [27:0] insn_o_1_97_0;
  wire  insn_o_1_98_0;
  wire  insn_o_1_99_0;
  wire  insn_o_1_100_0;
  wire  [0:0] insn_o_1_101_0;
  wire  [7:0] insn_o_1_102_0;
  wire  [27:0] insn_o_1_103_0;
  wire  [27:0] insn_o_1_104_0;
  wire  insn_o_1_105_0;
  wire  insn_o_1_106_0;
  wire  insn_o_1_107_0;
  wire  insn_o_1_108_0;
  wire  insn_o_1_109_0;
  wire  insn_o_1_110_0;
  wire  [27:0] insn_o_1_111_0;
  wire  [27:0] insn_o_1_112_0;
  wire  [27:0] insn_o_1_113_0;
  wire  [27:0] insn_o_1_114_0;
  wire  [27:0] insn_o_1_115_0;
  wire  insn_o_1_116_0;
  wire  insn_o_1_117_0;
  wire  [7:0] insn_o_1_118_0;
  wire  [0:0] insn_o_1_119_0;
  wire  insn_o_1_120_0;
  wire  insn_o_1_121_0;
  wire  insn_o_1_122_0;
  wire  insn_o_1_123_0;
  wire  insn_o_1_124_0;
  wire  insn_o_1_125_0;
  wire  [27:0] insn_o_1_126_0;
  wire  [15:0] insn_o_1_127_0;
  wire  [0:0] insn_o_1_128_0;
  wire  [11:0] insn_o_1_129_0;
  wire  [27:0] insn_o_1_130_0;
  wire  [27:0] insn_o_1_131_0;
  wire  [7:0] insn_o_1_132_0;
  wire  [0:0] insn_o_1_133_0;
  wire  [19:0] insn_o_1_134_0;
  wire  [27:0] insn_o_1_135_0;
  wire  [27:0] insn_o_1_136_0;
  wire  [3:0] insn_o_1_137_0;
  wire  [0:0] insn_o_1_138_0;
  wire  [23:0] insn_o_1_139_0;
  wire  [27:0] insn_o_1_140_0;
  wire  [27:0] insn_o_1_141_0;
  wire  [1:0] insn_o_1_142_0;
  wire  [0:0] insn_o_1_143_0;
  wire  [25:0] insn_o_1_144_0;
  wire  [27:0] insn_o_1_145_0;
  wire  [27:0] insn_o_1_146_0;
  wire  [0:0] insn_o_1_147_0;
  wire  [0:0] insn_o_1_148_0;
  wire  [26:0] insn_o_1_149_0;
  wire  [27:0] insn_o_1_150_0;
  wire  [27:0] insn_o_1_151_0;
  wire  [4:0] insn_o_1_152_0;
  wire  signed [8:0] insn_o_1_153_0;
  wire  signed [8:0] insn_o_1_154_0;
  wire  [27:0] insn_o_1_155_0;
  wire  [0:0] insn_o_1_156_0;
  wire  insn_o_1_157_0;
  wire  insn_o_1_158_0;
  wire  insn_o_1_159_0;
  wire  insn_o_1_160_0;
  wire  insn_o_1_161_0;
  wire  insn_o_1_162_0;
  wire  insn_o_1_163_0;
  wire  insn_o_1_164_0;
  wire  [23:0] insn_o_1_165_0;
  wire  [0:0] insn_o_1_166_0;
  wire  [0:0] insn_o_1_167_0;
  wire  [0:0] insn_o_1_168_0;
  wire  [0:0] insn_o_1_169_0;
  wire  [0:0] insn_o_1_170_0;
  wire  [0:0] insn_o_1_171_0;
  wire  [0:0] insn_o_1_172_0;
  wire  [0:0] insn_o_1_173_0;
  wire  [0:0] insn_o_1_174_0;
  wire  [23:0] insn_o_1_175_0;
  wire  insn_o_1_176_0;
  wire  [0:0] insn_o_1_177_0;
  wire  signed [8:0] insn_o_1_178_0;
  wire  [0:0] insn_o_1_179_0;
  wire  insn_o_1_180_0;
  wire  insn_o_1_181_0;
  wire  insn_o_1_182_0;
  wire  insn_o_1_183_0;
  wire  insn_o_1_184_0;
  wire  insn_o_1_185_0;
  wire  insn_o_1_186_0;
  wire  insn_o_1_187_0;
  wire  insn_o_1_188_0;
  wire  insn_o_1_189_0;
  wire  insn_o_1_190_0;
  wire  insn_o_1_191_0;
  wire  insn_o_1_192_0;
  wire  insn_o_1_193_0;
  wire  insn_o_1_194_0;
  wire  insn_o_1_195_0;
  wire  [0:0] insn_o_1_196_0;
  wire  [22:0] insn_o_1_197_0;
  wire  [7:0] insn_o_1_198_0;
  wire  insn_o_1_199_0;
  wire  insn_o_1_200_0;
  wire  [0:0] insn_o_1_201_0;
  wire  insn_o_1_202_0;
  wire  insn_o_1_203_0;
  wire  insn_o_1_204_0;
  wire  [0:0] insn_o_1_205_0;
  wire  [22:0] insn_o_1_206_0;
  wire  [7:0] insn_o_1_207_0;
  wire  [0:0] insn_o_1_208_0;
  wire  [22:0] insn_o_1_209_0;
  wire  [7:0] insn_o_1_210_0;
  wire  [0:0] insn_o_1_211_0;
  wire  [22:0] insn_o_1_212_0;
  wire  [7:0] insn_o_1_213_0;
  wire  [0:0] insn_o_1_214_0;
  wire  [22:0] insn_o_1_215_0;
  wire  [7:0] insn_o_1_216_0;
  wire  [0:0] insn_o_1_217_0;
  wire  [22:0] insn_o_1_218_0;
  wire  [7:0] insn_o_1_219_0;
  wire  [0:0] insn_o_1_220_0;
  wire  [31:0] insn_o_1_221_0;
  // Insn assigns
  assign insn_o_1_9_0 = i_valid;
  assign start = insn_o_1_9_0;
  assign insn_o_1_10_0 = sub;
  assign insn_o_1_11_0 = a_in;
  assign stage1_a_data_in = insn_o_1_11_0;
  assign insn_o_1_12_0 = stage1_a_data_in[22:0];
  assign stage1_a_fraction_in = insn_o_1_12_0;
  assign insn_o_1_13_0 = stage1_a_data_in[30:23];
  assign stage1_a_exponent_in = insn_o_1_13_0;
  assign insn_o_1_14_0 = stage1_a_data_in[31:31];
  assign insn_o_1_17_0 = b_in;
  assign stage1_b_data_in = insn_o_1_17_0;
  assign insn_o_1_18_0 = stage1_b_data_in[22:0];
  assign stage1_b_fraction_in = insn_o_1_18_0;
  assign insn_o_1_19_0 = stage1_b_data_in[30:23];
  assign stage1_b_exponent_in = insn_o_1_19_0;
  assign insn_o_1_20_0 = stage1_b_data_in[31:31];
  assign insn_o_1_23_0 = eq_18_d0;
  assign stage2_a_exponent_is_all_1 = insn_o_1_23_0;
  assign insn_o_1_24_0 = eq_19_d0;
  assign stage2_a_exponent_is_all_0 = insn_o_1_24_0;
  assign insn_o_1_25_0 = eq_20_d0;
  assign stage2_a_fraction_is_all_0 = insn_o_1_25_0;
  assign insn_o_1_26_0 = ~stage2_a_fraction_is_all_0;
  assign stage2_a_fraction_is_not_0 = insn_o_1_26_0;
  assign insn_o_1_27_0 = ~stage2_a_exponent_is_all_0;
  assign stage2_a_fraction_msb = insn_o_1_27_0;
  assign insn_o_1_28_0 = {stage2_a_fraction_msb, stage1_a_fraction};
  assign stage2_a_fraction_in = insn_o_1_28_0;
  assign stage2_a_exponent_in = stage1_a_exponent;
  assign stage2_a_sign_in = stage1_a_sign;
  assign insn_o_1_31_0 = stage2_a_exponent_is_all_0 & stage2_a_fraction_is_all_0;
  assign insn_o_1_32_0 = stage2_a_exponent_is_all_1 & stage2_a_fraction_is_all_0;
  assign insn_o_1_33_0 = stage2_a_exponent_is_all_1 & stage2_a_fraction_is_not_0;
  assign insn_o_1_34_0 = eq_29_d0;
  assign stage2_b_exponent_is_all_1 = insn_o_1_34_0;
  assign insn_o_1_35_0 = eq_30_d0;
  assign stage2_b_exponent_is_all_0 = insn_o_1_35_0;
  assign insn_o_1_36_0 = eq_31_d0;
  assign stage2_b_fraction_is_all_0 = insn_o_1_36_0;
  assign insn_o_1_37_0 = ~stage2_b_fraction_is_all_0;
  assign stage2_b_fraction_is_not_0 = insn_o_1_37_0;
  assign insn_o_1_38_0 = ~stage2_b_exponent_is_all_0;
  assign stage2_b_fraction_msb = insn_o_1_38_0;
  assign insn_o_1_39_0 = {stage2_b_fraction_msb, stage1_b_fraction};
  assign stage2_b_fraction_in = insn_o_1_39_0;
  assign stage2_b_exponent_in = stage1_b_exponent;
  assign stage2_b_sign_in = stage1_b_sign;
  assign insn_o_1_42_0 = stage2_b_exponent_is_all_0 & stage2_b_fraction_is_all_0;
  assign insn_o_1_43_0 = stage2_b_exponent_is_all_1 & stage2_b_fraction_is_all_0;
  assign insn_o_1_44_0 = stage2_b_exponent_is_all_1 & stage2_b_fraction_is_not_0;
  assign insn_o_1_45_0 = {stage1_a_exponent, stage1_a_fraction};
  assign stage2_a_abs_data = insn_o_1_45_0;
  assign insn_o_1_46_0 = {stage1_b_exponent, stage1_b_fraction};
  assign stage2_b_abs_data = insn_o_1_46_0;
  assign insn_o_1_47_0 = gt_42_d0;
  assign stage2_b_gt_a_125 = insn_o_1_47_0;
  assign insn_o_1_48_0 = stage2_b_gt_a_125 ? stage2_b_fraction_in : stage2_a_fraction_in;
  assign insn_o_1_49_0 = stage2_b_gt_a_125 ? stage2_b_exponent_in : stage2_a_exponent_in;
  assign insn_o_1_50_0 = stage2_b_gt_a_125 ? stage2_b_sign_in : stage2_a_sign_in;
  assign insn_o_1_51_0 = stage2_b_gt_a_125 ? stage2_a_fraction_in : stage2_b_fraction_in;
  assign insn_o_1_52_0 = stage2_b_gt_a_125 ? stage2_a_exponent_in : stage2_b_exponent_in;
  assign insn_o_1_53_0 = stage2_b_gt_a_125 ? stage2_a_sign_in : stage2_b_sign_in;
  assign insn_o_1_56_0 = stage2_sub ^ stage2_l_sign;
  assign stage3_sub_xor_l_sign = insn_o_1_56_0;
  assign insn_o_1_57_0 = stage2_b_gt_a ? stage3_sub_xor_l_sign : stage2_l_sign;
  assign insn_o_1_58_0 = stage2_s_sign ^ stage3_sub_xor_l_sign;
  assign insn_o_1_59_0 = sub_54_d0;
  assign insn_o_1_71_0 = {1'd0, stage3_s_fraction, 27'd0};
  assign stage4_shift_fractions_0 = insn_o_1_71_0;
  assign insn_o_1_72_0 = stage3_diff_exponent[0:0];
  assign anon_141 = insn_o_1_72_0;
  assign insn_o_1_73_0 = stage4_shift_fractions_0[51:1];
  assign anon_142 = insn_o_1_73_0;
  assign insn_o_1_74_0 = {1'd0, anon_142};
  assign anon_143 = insn_o_1_74_0;
  assign insn_o_1_75_0 = anon_141 ? anon_143 : stage4_shift_fractions_0;
  assign stage4_shift_fractions_1 = insn_o_1_75_0;
  assign insn_o_1_76_0 = stage3_diff_exponent[1:1];
  assign anon_149 = insn_o_1_76_0;
  assign insn_o_1_77_0 = stage4_shift_fractions_1[51:2];
  assign anon_150 = insn_o_1_77_0;
  assign insn_o_1_78_0 = {2'd0, anon_150};
  assign anon_151 = insn_o_1_78_0;
  assign insn_o_1_79_0 = anon_149 ? anon_151 : stage4_shift_fractions_1;
  assign stage4_shift_fractions_2 = insn_o_1_79_0;
  assign insn_o_1_80_0 = stage3_diff_exponent[2:2];
  assign anon_157 = insn_o_1_80_0;
  assign insn_o_1_81_0 = stage4_shift_fractions_2[51:4];
  assign anon_158 = insn_o_1_81_0;
  assign insn_o_1_82_0 = {4'd0, anon_158};
  assign anon_159 = insn_o_1_82_0;
  assign insn_o_1_83_0 = anon_157 ? anon_159 : stage4_shift_fractions_2;
  assign stage4_shift_fractions_3 = insn_o_1_83_0;
  assign insn_o_1_84_0 = stage3_diff_exponent[3:3];
  assign anon_165 = insn_o_1_84_0;
  assign insn_o_1_85_0 = stage4_shift_fractions_3[51:8];
  assign anon_166 = insn_o_1_85_0;
  assign insn_o_1_86_0 = {8'd0, anon_166};
  assign anon_167 = insn_o_1_86_0;
  assign insn_o_1_87_0 = anon_165 ? anon_167 : stage4_shift_fractions_3;
  assign stage4_shift_fractions_4 = insn_o_1_87_0;
  assign insn_o_1_88_0 = stage3_diff_exponent[4:4];
  assign anon_173 = insn_o_1_88_0;
  assign insn_o_1_89_0 = stage4_shift_fractions_4[51:16];
  assign anon_174 = insn_o_1_89_0;
  assign insn_o_1_90_0 = {16'd0, anon_174};
  assign anon_175 = insn_o_1_90_0;
  assign insn_o_1_91_0 = anon_173 ? anon_175 : stage4_shift_fractions_4;
  assign stage4_shift_fractions_5 = insn_o_1_91_0;
  assign insn_o_1_92_0 = gte_87_d0;
  assign stage4_s_under = insn_o_1_92_0;
  assign insn_o_1_93_0 = stage4_shift_fractions_5[51:25];
  assign stage4_s_fraction_data = insn_o_1_93_0;
  assign insn_o_1_94_0 = stage4_shift_fractions_5[24:0];
  assign stage4_s_sticky_data = insn_o_1_94_0;
  assign insn_o_1_95_0 = eq_90_d0;
  assign anon_191 = insn_o_1_95_0;
  assign insn_o_1_96_0 = ~anon_191;
  assign stage4_s_sticky = insn_o_1_96_0;
  assign insn_o_1_97_0 = {stage4_s_fraction_data, stage4_s_sticky};
  assign stage4_s_fraction_181 = insn_o_1_97_0;
  assign insn_o_1_103_0 = stage4_s_under ? 28'd1 : stage4_s_fraction_181;
  assign insn_o_1_104_0 = {1'd0, stage3_l_fraction, 3'd0};
  assign stage5_add_s_fraction = stage4_s_fraction;
  assign insn_o_1_112_0 = ~stage4_s_fraction;
  assign anon_196 = insn_o_1_112_0;
  assign insn_o_1_113_0 = add_108_d0;
  assign stage5_sub_s_fraction = insn_o_1_113_0;
  assign insn_o_1_114_0 = stage4_op_sub ? stage5_sub_s_fraction : stage5_add_s_fraction;
  assign stage5_s_fraction = insn_o_1_114_0;
  assign insn_o_1_115_0 = add_110_d0;
  assign stage6_fraction_data_5 = stage5_t_fraction;
  assign insn_o_1_127_0 = stage6_fraction_data_5[27:12];
  assign anon_214 = insn_o_1_127_0;
  assign insn_o_1_128_0 = eq_123_d0;
  assign stage6_shift_flag_4 = insn_o_1_128_0;
  assign insn_o_1_129_0 = stage6_fraction_data_5[11:0];
  assign anon_218 = insn_o_1_129_0;
  assign insn_o_1_130_0 = {anon_218, 16'd0};
  assign anon_219 = insn_o_1_130_0;
  assign insn_o_1_131_0 = stage6_shift_flag_4 ? anon_219 : stage6_fraction_data_5;
  assign stage6_fraction_data_4 = insn_o_1_131_0;
  assign insn_o_1_132_0 = stage6_fraction_data_4[27:20];
  assign anon_223 = insn_o_1_132_0;
  assign insn_o_1_133_0 = eq_128_d0;
  assign stage6_shift_flag_3 = insn_o_1_133_0;
  assign insn_o_1_134_0 = stage6_fraction_data_4[19:0];
  assign anon_227 = insn_o_1_134_0;
  assign insn_o_1_135_0 = {anon_227, 8'd0};
  assign anon_228 = insn_o_1_135_0;
  assign insn_o_1_136_0 = stage6_shift_flag_3 ? anon_228 : stage6_fraction_data_4;
  assign stage6_fraction_data_3 = insn_o_1_136_0;
  assign insn_o_1_137_0 = stage6_fraction_data_3[27:24];
  assign anon_232 = insn_o_1_137_0;
  assign insn_o_1_138_0 = eq_133_d0;
  assign stage6_shift_flag_2 = insn_o_1_138_0;
  assign insn_o_1_139_0 = stage6_fraction_data_3[23:0];
  assign anon_236 = insn_o_1_139_0;
  assign insn_o_1_140_0 = {anon_236, 4'd0};
  assign anon_237 = insn_o_1_140_0;
  assign insn_o_1_141_0 = stage6_shift_flag_2 ? anon_237 : stage6_fraction_data_3;
  assign stage6_fraction_data_2 = insn_o_1_141_0;
  assign insn_o_1_142_0 = stage6_fraction_data_2[27:26];
  assign anon_241 = insn_o_1_142_0;
  assign insn_o_1_143_0 = eq_138_d0;
  assign stage6_shift_flag_1 = insn_o_1_143_0;
  assign insn_o_1_144_0 = stage6_fraction_data_2[25:0];
  assign anon_245 = insn_o_1_144_0;
  assign insn_o_1_145_0 = {anon_245, 2'd0};
  assign anon_246 = insn_o_1_145_0;
  assign insn_o_1_146_0 = stage6_shift_flag_1 ? anon_246 : stage6_fraction_data_2;
  assign stage6_fraction_data_1 = insn_o_1_146_0;
  assign insn_o_1_147_0 = stage6_fraction_data_1[27:27];
  assign anon_250 = insn_o_1_147_0;
  assign insn_o_1_148_0 = eq_143_d0;
  assign stage6_shift_flag_0 = insn_o_1_148_0;
  assign insn_o_1_149_0 = stage6_fraction_data_1[26:0];
  assign anon_254 = insn_o_1_149_0;
  assign insn_o_1_150_0 = {anon_254, 1'd0};
  assign anon_255 = insn_o_1_150_0;
  assign insn_o_1_151_0 = stage6_shift_flag_0 ? anon_255 : stage6_fraction_data_1;
  assign stage6_fraction_data_0 = insn_o_1_151_0;
  assign insn_o_1_152_0 = {stage6_shift_flag_4, stage6_shift_flag_3, stage6_shift_flag_2, stage6_shift_flag_1, stage6_shift_flag_0};
  assign stage6_shift = insn_o_1_152_0;
  assign insn_o_1_153_0 = sub_148_d0;
  assign anon_257 = insn_o_1_153_0;
  assign insn_o_1_154_0 = add_149_d0;
  assign insn_o_1_165_0 = stage6_t_fraction[27:4];
  assign stage7_fraction_data = insn_o_1_165_0;
  assign insn_o_1_166_0 = stage6_t_fraction[4:4];
  assign stage7_ulp = insn_o_1_166_0;
  assign insn_o_1_167_0 = stage6_t_fraction[3:3];
  assign stage7_uulp1 = insn_o_1_167_0;
  assign insn_o_1_168_0 = stage6_t_fraction[2:2];
  assign stage7_uulp2 = insn_o_1_168_0;
  assign insn_o_1_169_0 = stage6_t_fraction[1:1];
  assign stage7_uulp3 = insn_o_1_169_0;
  assign insn_o_1_170_0 = stage6_t_fraction[0:0];
  assign stage7_uulp4 = insn_o_1_170_0;
  assign insn_o_1_171_0 = stage7_ulp | stage7_uulp2;
  assign anon_278 = insn_o_1_171_0;
  assign insn_o_1_172_0 = anon_278 | stage7_uulp3;
  assign anon_279 = insn_o_1_172_0;
  assign insn_o_1_173_0 = anon_279 | stage7_uulp4;
  assign anon_280 = insn_o_1_173_0;
  assign insn_o_1_174_0 = stage7_uulp1 & anon_280;
  assign stage7_increment = insn_o_1_174_0;
  assign insn_o_1_175_0 = add_170_d0;
  assign insn_o_1_176_0 = eq_171_d0;
  assign anon_281 = insn_o_1_176_0;
  assign insn_o_1_177_0 = stage7_increment & anon_281;
  assign anon_282 = insn_o_1_177_0;
  assign insn_o_1_178_0 = add_173_d0;
  assign insn_o_1_188_0 = stage7_a_is_nan | stage7_b_is_nan;
  assign anon_293 = insn_o_1_188_0;
  assign insn_o_1_189_0 = stage7_a_is_inf & stage7_b_is_inf;
  assign anon_294 = insn_o_1_189_0;
  assign insn_o_1_190_0 = anon_294 & stage7_sub;
  assign anon_295 = insn_o_1_190_0;
  assign insn_o_1_191_0 = anon_293 | anon_295;
  assign stage8_set_nan = insn_o_1_191_0;
  assign insn_o_1_192_0 = ~stage8_set_nan;
  assign anon_296 = insn_o_1_192_0;
  assign insn_o_1_193_0 = stage7_a_is_inf | stage7_b_is_inf;
  assign anon_297 = insn_o_1_193_0;
  assign insn_o_1_194_0 = anon_296 & anon_297;
  assign stage8_set_inf = insn_o_1_194_0;
  assign insn_o_1_195_0 = stage7_a_is_zero & stage7_b_is_zero;
  assign stage8_set_zero = insn_o_1_195_0;
  assign insn_o_1_196_0 = stage7_t_fraction[23:23];
  assign stage8_fraction_msb = insn_o_1_196_0;
  assign insn_o_1_197_0 = stage7_t_fraction[22:0];
  assign stage8_fraction_in = insn_o_1_197_0;
  assign insn_o_1_198_0 = stage7_t_exponent[7:0];
  assign stage8_exponent_in = insn_o_1_198_0;
  assign insn_o_1_199_0 = gt_194_d0;
  assign stage8_exp_natural = insn_o_1_199_0;
  assign insn_o_1_200_0 = ~stage8_exp_natural;
  assign anon_312 = insn_o_1_200_0;
  assign insn_o_1_201_0 = ~stage8_fraction_msb;
  assign anon_313 = insn_o_1_201_0;
  assign insn_o_1_202_0 = anon_312 | anon_313;
  assign stage8_exp_underflow = insn_o_1_202_0;
  assign insn_o_1_203_0 = gte_198_d0;
  assign anon_315 = insn_o_1_203_0;
  assign insn_o_1_204_0 = anon_315 & stage8_fraction_msb;
  assign stage8_exp_overflow = insn_o_1_204_0;
  assign stage8_sign_in = stage7_t_sign;
  assign insn_o_1_206_0 = stage8_exp_overflow ? 23'd0 : stage8_fraction_in;
  assign stage8_fraction_i1 = insn_o_1_206_0;
  assign insn_o_1_207_0 = stage8_exp_overflow ? 8'd255 : stage8_exponent_in;
  assign stage8_exponent_i1 = insn_o_1_207_0;
  assign stage8_sign_i1 = stage8_sign_in;
  assign insn_o_1_209_0 = stage8_exp_underflow ? 23'd0 : stage8_fraction_i1;
  assign stage8_fraction_i2 = insn_o_1_209_0;
  assign insn_o_1_210_0 = stage8_exp_underflow ? 8'd0 : stage8_exponent_i1;
  assign stage8_exponent_i2 = insn_o_1_210_0;
  assign stage8_sign_i2 = stage8_sign_i1;
  assign insn_o_1_212_0 = stage8_set_nan ? 23'd2097152 : stage8_fraction_i2;
  assign stage8_fraction_i3 = insn_o_1_212_0;
  assign insn_o_1_213_0 = stage8_set_nan ? 8'd255 : stage8_exponent_i2;
  assign stage8_exponent_i3 = insn_o_1_213_0;
  assign insn_o_1_214_0 = stage8_set_nan ? 1'd0 : stage8_sign_i2;
  assign stage8_sign_i3 = insn_o_1_214_0;
  assign insn_o_1_215_0 = stage8_set_inf ? 23'd0 : stage8_fraction_i3;
  assign stage8_fraction_i4 = insn_o_1_215_0;
  assign insn_o_1_216_0 = stage8_set_inf ? 8'd255 : stage8_exponent_i3;
  assign stage8_exponent_i4 = insn_o_1_216_0;
  assign stage8_sign_i4 = stage8_sign_i3;
  assign insn_o_1_218_0 = stage8_set_zero ? 23'd0 : stage8_fraction_i4;
  assign stage8_fraction_o = insn_o_1_218_0;
  assign insn_o_1_219_0 = stage8_set_zero ? 8'd0 : stage8_exponent_i4;
  assign stage8_exponent_o = insn_o_1_219_0;
  assign stage8_sign_o = stage8_sign_i4;
  assign insn_o_1_221_0 = {stage8_sign_o, stage8_exponent_o, stage8_fraction_o};
  assign stage8_result = insn_o_1_221_0;

  // Table 1
  always @(posedge clk) begin
    if (!rst_n) begin
      st_1_1 <= 0;
      st_1_2 <= 0;
      st_1_3 <= 0;
      st_1_4 <= 0;
      st_1_5 <= 0;
      st_1_6 <= 0;
      st_1_7 <= 0;
      st_1_8 <= 0;
    end else begin
      if (start) begin
          stage1_a_fraction <= stage1_a_fraction_in;
          stage1_a_exponent <= stage1_a_exponent_in;
          stage1_b_fraction <= stage1_b_fraction_in;
          stage1_b_exponent <= stage1_b_exponent_in;
          stage1_sub <= insn_o_1_10_0;
          stage1_a_sign <= insn_o_1_14_0;
          stage1_b_sign <= insn_o_1_20_0;
      end
      st_1_2 <= start;
      if (st_1_2) begin
          stage2_b_gt_a <= stage2_b_gt_a_125;
          stage2_sub <= stage1_sub;
          stage2_a_is_zero <= insn_o_1_31_0;
          stage2_a_is_inf <= insn_o_1_32_0;
          stage2_a_is_nan <= insn_o_1_33_0;
          stage2_b_is_zero <= insn_o_1_42_0;
          stage2_b_is_inf <= insn_o_1_43_0;
          stage2_b_is_nan <= insn_o_1_44_0;
          stage2_l_fraction <= insn_o_1_48_0;
          stage2_l_exponent <= insn_o_1_49_0;
          stage2_l_sign <= insn_o_1_50_0;
          stage2_s_fraction <= insn_o_1_51_0;
          stage2_s_exponent <= insn_o_1_52_0;
          stage2_s_sign <= insn_o_1_53_0;
      end
      st_1_3 <= st_1_2;
      if (st_1_3) begin
          stage3_t_exponent <= stage2_l_exponent;
          stage3_l_fraction <= stage2_l_fraction;
          stage3_s_fraction <= stage2_s_fraction;
          stage3_b_gt_a <= stage2_b_gt_a;
          stage3_sub <= stage2_sub;
          stage3_a_is_zero <= stage2_a_is_zero;
          stage3_a_is_inf <= stage2_a_is_inf;
          stage3_a_is_nan <= stage2_a_is_nan;
          stage3_b_is_zero <= stage2_b_is_zero;
          stage3_b_is_inf <= stage2_b_is_inf;
          stage3_b_is_nan <= stage2_b_is_nan;
          stage3_t_sign <= insn_o_1_57_0;
          stage3_op_sub <= insn_o_1_58_0;
          stage3_diff_exponent <= insn_o_1_59_0;
      end
      st_1_4 <= st_1_3;
      if (st_1_4) begin
          stage4_sub <= stage3_sub;
          stage4_op_sub <= stage3_op_sub;
          stage4_b_gt_a <= stage3_b_gt_a;
          stage4_t_sign <= stage3_t_sign;
          stage4_t_exponent <= stage3_t_exponent;
          stage4_a_is_zero <= stage3_a_is_zero;
          stage4_a_is_inf <= stage3_a_is_inf;
          stage4_a_is_nan <= stage3_a_is_nan;
          stage4_b_is_zero <= stage3_b_is_zero;
          stage4_b_is_inf <= stage3_b_is_inf;
          stage4_b_is_nan <= stage3_b_is_nan;
          stage4_s_fraction <= insn_o_1_103_0;
          stage4_l_fraction <= insn_o_1_104_0;
      end
      st_1_5 <= st_1_4;
      if (st_1_5) begin
          stage5_sub <= stage4_sub;
          stage5_b_gt_a <= stage4_b_gt_a;
          stage5_t_exponent <= stage4_t_exponent;
          stage5_t_sign <= stage4_t_sign;
          stage5_a_is_zero <= stage4_a_is_zero;
          stage5_a_is_inf <= stage4_a_is_inf;
          stage5_a_is_nan <= stage4_a_is_nan;
          stage5_b_is_zero <= stage4_b_is_zero;
          stage5_b_is_inf <= stage4_b_is_inf;
          stage5_b_is_nan <= stage4_b_is_nan;
          stage5_t_fraction <= insn_o_1_115_0;
      end
      st_1_6 <= st_1_5;
      if (st_1_6) begin
          stage6_t_fraction <= stage6_fraction_data_0;
          stage6_t_sign <= stage5_t_sign;
          stage6_sub <= stage5_sub;
          stage6_b_gt_a <= stage5_b_gt_a;
          stage6_a_is_zero <= stage5_a_is_zero;
          stage6_a_is_inf <= stage5_a_is_inf;
          stage6_a_is_nan <= stage5_a_is_nan;
          stage6_b_is_zero <= stage5_b_is_zero;
          stage6_b_is_inf <= stage5_b_is_inf;
          stage6_b_is_nan <= stage5_b_is_nan;
          stage6_t_exponent <= insn_o_1_154_0;
      end
      st_1_7 <= st_1_6;
      if (st_1_7) begin
          stage7_t_sign <= stage6_t_sign;
          stage7_sub <= stage6_sub;
          stage7_b_gt_a <= stage6_b_gt_a;
          stage7_a_is_zero <= stage6_a_is_zero;
          stage7_a_is_inf <= stage6_a_is_inf;
          stage7_a_is_nan <= stage6_a_is_nan;
          stage7_b_is_zero <= stage6_b_is_zero;
          stage7_b_is_inf <= stage6_b_is_inf;
          stage7_b_is_nan <= stage6_b_is_nan;
          stage7_t_fraction <= insn_o_1_175_0;
          stage7_t_exponent <= insn_o_1_178_0;
      end
      st_1_8 <= st_1_7;
      if (st_1_8) begin
          z_out <= stage8_result;
      end
    end
  end

endmodule
