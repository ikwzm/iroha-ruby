// Generated from iroha-0.1.0.

module div(clk, rst_n, i_valid, dividend, divisor, quotient, remainder, o_valid);
  input clk;
  input rst_n;
  input i_valid;
  input [31:0] dividend;
  input [15:0] divisor;
  output [31:0] quotient;
  output [15:0] remainder;
  output o_valid;
  reg [31:0] quotient;
  reg [15:0] remainder;
  reg o_valid;

  // State decls
  reg st_1_1;
  reg st_1_2;
  reg st_1_3;
  reg st_1_4;
  reg st_1_5;
  reg st_1_6;
  reg st_1_7;
  reg st_1_8;
  reg st_1_9;
  reg st_1_10;
  reg st_1_11;
  reg st_1_12;
  reg st_1_13;
  reg st_1_14;
  reg st_1_15;
  reg st_1_16;
  reg st_1_17;
  reg st_1_18;
  reg st_1_19;
  reg st_1_20;
  reg st_1_21;
  reg st_1_22;
  reg st_1_23;
  reg st_1_24;
  reg st_1_25;
  reg st_1_26;
  reg st_1_27;
  reg st_1_28;
  reg st_1_29;
  reg st_1_30;
  reg st_1_31;
  reg st_1_32;
  reg st_1_33;
  // State vars
  // Registers
  wire  [0:0] start;
  reg  [47:0] zi_00;
  reg  [47:0] zi_01;
  reg  [47:0] zi_02;
  reg  [47:0] zi_03;
  reg  [47:0] zi_04;
  reg  [47:0] zi_05;
  reg  [47:0] zi_06;
  reg  [47:0] zi_07;
  reg  [47:0] zi_08;
  reg  [47:0] zi_09;
  reg  [47:0] zi_10;
  reg  [47:0] zi_11;
  reg  [47:0] zi_12;
  reg  [47:0] zi_13;
  reg  [47:0] zi_14;
  reg  [47:0] zi_15;
  reg  [47:0] zi_16;
  reg  [47:0] zi_17;
  reg  [47:0] zi_18;
  reg  [47:0] zi_19;
  reg  [47:0] zi_20;
  reg  [47:0] zi_21;
  reg  [47:0] zi_22;
  reg  [47:0] zi_23;
  reg  [47:0] zi_24;
  reg  [47:0] zi_25;
  reg  [47:0] zi_26;
  reg  [47:0] zi_27;
  reg  [47:0] zi_28;
  reg  [47:0] zi_29;
  reg  [47:0] zi_30;
  reg  [47:0] zi_31;
  reg  [15:0] di_00;
  reg  [15:0] di_01;
  reg  [15:0] di_02;
  reg  [15:0] di_03;
  reg  [15:0] di_04;
  reg  [15:0] di_05;
  reg  [15:0] di_06;
  reg  [15:0] di_07;
  reg  [15:0] di_08;
  reg  [15:0] di_09;
  reg  [15:0] di_10;
  reg  [15:0] di_11;
  reg  [15:0] di_12;
  reg  [15:0] di_13;
  reg  [15:0] di_14;
  reg  [15:0] di_15;
  reg  [15:0] di_16;
  reg  [15:0] di_17;
  reg  [15:0] di_18;
  reg  [15:0] di_19;
  reg  [15:0] di_20;
  reg  [15:0] di_21;
  reg  [15:0] di_22;
  reg  [15:0] di_23;
  reg  [15:0] di_24;
  reg  [15:0] di_25;
  reg  [15:0] di_26;
  reg  [15:0] di_27;
  reg  [15:0] di_28;
  reg  [15:0] di_29;
  reg  [15:0] di_30;
  reg  [15:0] di_31;
  wire  [31:0] stage_32_zi_l;
  wire  [47:0] stage_32_zi_i;
  wire  [16:0] stage_31_pr;
  wire  [16:0] stage_31_sb;
  wire  [15:0] stage_31_m0;
  wire  [15:0] stage_31_m1;
  wire  [0:0] stage_31_ms;
  wire  [15:0] stage_31_mx;
  wire  [30:0] stage_31_zl;
  wire  [0:0] stage_31_zb;
  wire  [47:0] stage_31_zo;
  wire  [16:0] stage_30_pr;
  wire  [16:0] stage_30_sb;
  wire  [15:0] stage_30_m0;
  wire  [15:0] stage_30_m1;
  wire  [0:0] stage_30_ms;
  wire  [15:0] stage_30_mx;
  wire  [30:0] stage_30_zl;
  wire  [0:0] stage_30_zb;
  wire  [47:0] stage_30_zo;
  wire  [16:0] stage_29_pr;
  wire  [16:0] stage_29_sb;
  wire  [15:0] stage_29_m0;
  wire  [15:0] stage_29_m1;
  wire  [0:0] stage_29_ms;
  wire  [15:0] stage_29_mx;
  wire  [30:0] stage_29_zl;
  wire  [0:0] stage_29_zb;
  wire  [47:0] stage_29_zo;
  wire  [16:0] stage_28_pr;
  wire  [16:0] stage_28_sb;
  wire  [15:0] stage_28_m0;
  wire  [15:0] stage_28_m1;
  wire  [0:0] stage_28_ms;
  wire  [15:0] stage_28_mx;
  wire  [30:0] stage_28_zl;
  wire  [0:0] stage_28_zb;
  wire  [47:0] stage_28_zo;
  wire  [16:0] stage_27_pr;
  wire  [16:0] stage_27_sb;
  wire  [15:0] stage_27_m0;
  wire  [15:0] stage_27_m1;
  wire  [0:0] stage_27_ms;
  wire  [15:0] stage_27_mx;
  wire  [30:0] stage_27_zl;
  wire  [0:0] stage_27_zb;
  wire  [47:0] stage_27_zo;
  wire  [16:0] stage_26_pr;
  wire  [16:0] stage_26_sb;
  wire  [15:0] stage_26_m0;
  wire  [15:0] stage_26_m1;
  wire  [0:0] stage_26_ms;
  wire  [15:0] stage_26_mx;
  wire  [30:0] stage_26_zl;
  wire  [0:0] stage_26_zb;
  wire  [47:0] stage_26_zo;
  wire  [16:0] stage_25_pr;
  wire  [16:0] stage_25_sb;
  wire  [15:0] stage_25_m0;
  wire  [15:0] stage_25_m1;
  wire  [0:0] stage_25_ms;
  wire  [15:0] stage_25_mx;
  wire  [30:0] stage_25_zl;
  wire  [0:0] stage_25_zb;
  wire  [47:0] stage_25_zo;
  wire  [16:0] stage_24_pr;
  wire  [16:0] stage_24_sb;
  wire  [15:0] stage_24_m0;
  wire  [15:0] stage_24_m1;
  wire  [0:0] stage_24_ms;
  wire  [15:0] stage_24_mx;
  wire  [30:0] stage_24_zl;
  wire  [0:0] stage_24_zb;
  wire  [47:0] stage_24_zo;
  wire  [16:0] stage_23_pr;
  wire  [16:0] stage_23_sb;
  wire  [15:0] stage_23_m0;
  wire  [15:0] stage_23_m1;
  wire  [0:0] stage_23_ms;
  wire  [15:0] stage_23_mx;
  wire  [30:0] stage_23_zl;
  wire  [0:0] stage_23_zb;
  wire  [47:0] stage_23_zo;
  wire  [16:0] stage_22_pr;
  wire  [16:0] stage_22_sb;
  wire  [15:0] stage_22_m0;
  wire  [15:0] stage_22_m1;
  wire  [0:0] stage_22_ms;
  wire  [15:0] stage_22_mx;
  wire  [30:0] stage_22_zl;
  wire  [0:0] stage_22_zb;
  wire  [47:0] stage_22_zo;
  wire  [16:0] stage_21_pr;
  wire  [16:0] stage_21_sb;
  wire  [15:0] stage_21_m0;
  wire  [15:0] stage_21_m1;
  wire  [0:0] stage_21_ms;
  wire  [15:0] stage_21_mx;
  wire  [30:0] stage_21_zl;
  wire  [0:0] stage_21_zb;
  wire  [47:0] stage_21_zo;
  wire  [16:0] stage_20_pr;
  wire  [16:0] stage_20_sb;
  wire  [15:0] stage_20_m0;
  wire  [15:0] stage_20_m1;
  wire  [0:0] stage_20_ms;
  wire  [15:0] stage_20_mx;
  wire  [30:0] stage_20_zl;
  wire  [0:0] stage_20_zb;
  wire  [47:0] stage_20_zo;
  wire  [16:0] stage_19_pr;
  wire  [16:0] stage_19_sb;
  wire  [15:0] stage_19_m0;
  wire  [15:0] stage_19_m1;
  wire  [0:0] stage_19_ms;
  wire  [15:0] stage_19_mx;
  wire  [30:0] stage_19_zl;
  wire  [0:0] stage_19_zb;
  wire  [47:0] stage_19_zo;
  wire  [16:0] stage_18_pr;
  wire  [16:0] stage_18_sb;
  wire  [15:0] stage_18_m0;
  wire  [15:0] stage_18_m1;
  wire  [0:0] stage_18_ms;
  wire  [15:0] stage_18_mx;
  wire  [30:0] stage_18_zl;
  wire  [0:0] stage_18_zb;
  wire  [47:0] stage_18_zo;
  wire  [16:0] stage_17_pr;
  wire  [16:0] stage_17_sb;
  wire  [15:0] stage_17_m0;
  wire  [15:0] stage_17_m1;
  wire  [0:0] stage_17_ms;
  wire  [15:0] stage_17_mx;
  wire  [30:0] stage_17_zl;
  wire  [0:0] stage_17_zb;
  wire  [47:0] stage_17_zo;
  wire  [16:0] stage_16_pr;
  wire  [16:0] stage_16_sb;
  wire  [15:0] stage_16_m0;
  wire  [15:0] stage_16_m1;
  wire  [0:0] stage_16_ms;
  wire  [15:0] stage_16_mx;
  wire  [30:0] stage_16_zl;
  wire  [0:0] stage_16_zb;
  wire  [47:0] stage_16_zo;
  wire  [16:0] stage_15_pr;
  wire  [16:0] stage_15_sb;
  wire  [15:0] stage_15_m0;
  wire  [15:0] stage_15_m1;
  wire  [0:0] stage_15_ms;
  wire  [15:0] stage_15_mx;
  wire  [30:0] stage_15_zl;
  wire  [0:0] stage_15_zb;
  wire  [47:0] stage_15_zo;
  wire  [16:0] stage_14_pr;
  wire  [16:0] stage_14_sb;
  wire  [15:0] stage_14_m0;
  wire  [15:0] stage_14_m1;
  wire  [0:0] stage_14_ms;
  wire  [15:0] stage_14_mx;
  wire  [30:0] stage_14_zl;
  wire  [0:0] stage_14_zb;
  wire  [47:0] stage_14_zo;
  wire  [16:0] stage_13_pr;
  wire  [16:0] stage_13_sb;
  wire  [15:0] stage_13_m0;
  wire  [15:0] stage_13_m1;
  wire  [0:0] stage_13_ms;
  wire  [15:0] stage_13_mx;
  wire  [30:0] stage_13_zl;
  wire  [0:0] stage_13_zb;
  wire  [47:0] stage_13_zo;
  wire  [16:0] stage_12_pr;
  wire  [16:0] stage_12_sb;
  wire  [15:0] stage_12_m0;
  wire  [15:0] stage_12_m1;
  wire  [0:0] stage_12_ms;
  wire  [15:0] stage_12_mx;
  wire  [30:0] stage_12_zl;
  wire  [0:0] stage_12_zb;
  wire  [47:0] stage_12_zo;
  wire  [16:0] stage_11_pr;
  wire  [16:0] stage_11_sb;
  wire  [15:0] stage_11_m0;
  wire  [15:0] stage_11_m1;
  wire  [0:0] stage_11_ms;
  wire  [15:0] stage_11_mx;
  wire  [30:0] stage_11_zl;
  wire  [0:0] stage_11_zb;
  wire  [47:0] stage_11_zo;
  wire  [16:0] stage_10_pr;
  wire  [16:0] stage_10_sb;
  wire  [15:0] stage_10_m0;
  wire  [15:0] stage_10_m1;
  wire  [0:0] stage_10_ms;
  wire  [15:0] stage_10_mx;
  wire  [30:0] stage_10_zl;
  wire  [0:0] stage_10_zb;
  wire  [47:0] stage_10_zo;
  wire  [16:0] stage_9_pr;
  wire  [16:0] stage_9_sb;
  wire  [15:0] stage_9_m0;
  wire  [15:0] stage_9_m1;
  wire  [0:0] stage_9_ms;
  wire  [15:0] stage_9_mx;
  wire  [30:0] stage_9_zl;
  wire  [0:0] stage_9_zb;
  wire  [47:0] stage_9_zo;
  wire  [16:0] stage_8_pr;
  wire  [16:0] stage_8_sb;
  wire  [15:0] stage_8_m0;
  wire  [15:0] stage_8_m1;
  wire  [0:0] stage_8_ms;
  wire  [15:0] stage_8_mx;
  wire  [30:0] stage_8_zl;
  wire  [0:0] stage_8_zb;
  wire  [47:0] stage_8_zo;
  wire  [16:0] stage_7_pr;
  wire  [16:0] stage_7_sb;
  wire  [15:0] stage_7_m0;
  wire  [15:0] stage_7_m1;
  wire  [0:0] stage_7_ms;
  wire  [15:0] stage_7_mx;
  wire  [30:0] stage_7_zl;
  wire  [0:0] stage_7_zb;
  wire  [47:0] stage_7_zo;
  wire  [16:0] stage_6_pr;
  wire  [16:0] stage_6_sb;
  wire  [15:0] stage_6_m0;
  wire  [15:0] stage_6_m1;
  wire  [0:0] stage_6_ms;
  wire  [15:0] stage_6_mx;
  wire  [30:0] stage_6_zl;
  wire  [0:0] stage_6_zb;
  wire  [47:0] stage_6_zo;
  wire  [16:0] stage_5_pr;
  wire  [16:0] stage_5_sb;
  wire  [15:0] stage_5_m0;
  wire  [15:0] stage_5_m1;
  wire  [0:0] stage_5_ms;
  wire  [15:0] stage_5_mx;
  wire  [30:0] stage_5_zl;
  wire  [0:0] stage_5_zb;
  wire  [47:0] stage_5_zo;
  wire  [16:0] stage_4_pr;
  wire  [16:0] stage_4_sb;
  wire  [15:0] stage_4_m0;
  wire  [15:0] stage_4_m1;
  wire  [0:0] stage_4_ms;
  wire  [15:0] stage_4_mx;
  wire  [30:0] stage_4_zl;
  wire  [0:0] stage_4_zb;
  wire  [47:0] stage_4_zo;
  wire  [16:0] stage_3_pr;
  wire  [16:0] stage_3_sb;
  wire  [15:0] stage_3_m0;
  wire  [15:0] stage_3_m1;
  wire  [0:0] stage_3_ms;
  wire  [15:0] stage_3_mx;
  wire  [30:0] stage_3_zl;
  wire  [0:0] stage_3_zb;
  wire  [47:0] stage_3_zo;
  wire  [16:0] stage_2_pr;
  wire  [16:0] stage_2_sb;
  wire  [15:0] stage_2_m0;
  wire  [15:0] stage_2_m1;
  wire  [0:0] stage_2_ms;
  wire  [15:0] stage_2_mx;
  wire  [30:0] stage_2_zl;
  wire  [0:0] stage_2_zb;
  wire  [47:0] stage_2_zo;
  wire  [16:0] stage_1_pr;
  wire  [16:0] stage_1_sb;
  wire  [15:0] stage_1_m0;
  wire  [15:0] stage_1_m1;
  wire  [0:0] stage_1_ms;
  wire  [15:0] stage_1_mx;
  wire  [30:0] stage_1_zl;
  wire  [0:0] stage_1_zb;
  wire  [47:0] stage_1_zo;
  wire  [16:0] stage_0_pr;
  wire  [16:0] stage_0_sb;
  wire  [15:0] stage_0_m0;
  wire  [15:0] stage_0_m1;
  wire  [0:0] stage_0_ms;
  wire  [15:0] stage_0_mx;
  wire  [30:0] stage_0_zl;
  wire  [0:0] stage_0_zb;
  wire  [47:0] stage_0_zo;
  wire  [15:0] stage_0_zr;
  wire  [31:0] stage_0_zq;
  // Resources
  // sub:12
  wire [16:0] sub_12_s0;
  assign sub_12_s0 = stage_31_pr;
  wire [15:0] sub_12_s1;
  assign sub_12_s1 = di_31;
  wire [16:0] sub_12_d0;
  assign sub_12_d0 = sub_12_s0 - sub_12_s1;
  // sub:23
  wire [16:0] sub_23_s0;
  assign sub_23_s0 = stage_30_pr;
  wire [15:0] sub_23_s1;
  assign sub_23_s1 = di_30;
  wire [16:0] sub_23_d0;
  assign sub_23_d0 = sub_23_s0 - sub_23_s1;
  // sub:34
  wire [16:0] sub_34_s0;
  assign sub_34_s0 = stage_29_pr;
  wire [15:0] sub_34_s1;
  assign sub_34_s1 = di_29;
  wire [16:0] sub_34_d0;
  assign sub_34_d0 = sub_34_s0 - sub_34_s1;
  // sub:45
  wire [16:0] sub_45_s0;
  assign sub_45_s0 = stage_28_pr;
  wire [15:0] sub_45_s1;
  assign sub_45_s1 = di_28;
  wire [16:0] sub_45_d0;
  assign sub_45_d0 = sub_45_s0 - sub_45_s1;
  // sub:56
  wire [16:0] sub_56_s0;
  assign sub_56_s0 = stage_27_pr;
  wire [15:0] sub_56_s1;
  assign sub_56_s1 = di_27;
  wire [16:0] sub_56_d0;
  assign sub_56_d0 = sub_56_s0 - sub_56_s1;
  // sub:67
  wire [16:0] sub_67_s0;
  assign sub_67_s0 = stage_26_pr;
  wire [15:0] sub_67_s1;
  assign sub_67_s1 = di_26;
  wire [16:0] sub_67_d0;
  assign sub_67_d0 = sub_67_s0 - sub_67_s1;
  // sub:78
  wire [16:0] sub_78_s0;
  assign sub_78_s0 = stage_25_pr;
  wire [15:0] sub_78_s1;
  assign sub_78_s1 = di_25;
  wire [16:0] sub_78_d0;
  assign sub_78_d0 = sub_78_s0 - sub_78_s1;
  // sub:89
  wire [16:0] sub_89_s0;
  assign sub_89_s0 = stage_24_pr;
  wire [15:0] sub_89_s1;
  assign sub_89_s1 = di_24;
  wire [16:0] sub_89_d0;
  assign sub_89_d0 = sub_89_s0 - sub_89_s1;
  // sub:100
  wire [16:0] sub_100_s0;
  assign sub_100_s0 = stage_23_pr;
  wire [15:0] sub_100_s1;
  assign sub_100_s1 = di_23;
  wire [16:0] sub_100_d0;
  assign sub_100_d0 = sub_100_s0 - sub_100_s1;
  // sub:111
  wire [16:0] sub_111_s0;
  assign sub_111_s0 = stage_22_pr;
  wire [15:0] sub_111_s1;
  assign sub_111_s1 = di_22;
  wire [16:0] sub_111_d0;
  assign sub_111_d0 = sub_111_s0 - sub_111_s1;
  // sub:122
  wire [16:0] sub_122_s0;
  assign sub_122_s0 = stage_21_pr;
  wire [15:0] sub_122_s1;
  assign sub_122_s1 = di_21;
  wire [16:0] sub_122_d0;
  assign sub_122_d0 = sub_122_s0 - sub_122_s1;
  // sub:133
  wire [16:0] sub_133_s0;
  assign sub_133_s0 = stage_20_pr;
  wire [15:0] sub_133_s1;
  assign sub_133_s1 = di_20;
  wire [16:0] sub_133_d0;
  assign sub_133_d0 = sub_133_s0 - sub_133_s1;
  // sub:144
  wire [16:0] sub_144_s0;
  assign sub_144_s0 = stage_19_pr;
  wire [15:0] sub_144_s1;
  assign sub_144_s1 = di_19;
  wire [16:0] sub_144_d0;
  assign sub_144_d0 = sub_144_s0 - sub_144_s1;
  // sub:155
  wire [16:0] sub_155_s0;
  assign sub_155_s0 = stage_18_pr;
  wire [15:0] sub_155_s1;
  assign sub_155_s1 = di_18;
  wire [16:0] sub_155_d0;
  assign sub_155_d0 = sub_155_s0 - sub_155_s1;
  // sub:166
  wire [16:0] sub_166_s0;
  assign sub_166_s0 = stage_17_pr;
  wire [15:0] sub_166_s1;
  assign sub_166_s1 = di_17;
  wire [16:0] sub_166_d0;
  assign sub_166_d0 = sub_166_s0 - sub_166_s1;
  // sub:177
  wire [16:0] sub_177_s0;
  assign sub_177_s0 = stage_16_pr;
  wire [15:0] sub_177_s1;
  assign sub_177_s1 = di_16;
  wire [16:0] sub_177_d0;
  assign sub_177_d0 = sub_177_s0 - sub_177_s1;
  // sub:188
  wire [16:0] sub_188_s0;
  assign sub_188_s0 = stage_15_pr;
  wire [15:0] sub_188_s1;
  assign sub_188_s1 = di_15;
  wire [16:0] sub_188_d0;
  assign sub_188_d0 = sub_188_s0 - sub_188_s1;
  // sub:199
  wire [16:0] sub_199_s0;
  assign sub_199_s0 = stage_14_pr;
  wire [15:0] sub_199_s1;
  assign sub_199_s1 = di_14;
  wire [16:0] sub_199_d0;
  assign sub_199_d0 = sub_199_s0 - sub_199_s1;
  // sub:210
  wire [16:0] sub_210_s0;
  assign sub_210_s0 = stage_13_pr;
  wire [15:0] sub_210_s1;
  assign sub_210_s1 = di_13;
  wire [16:0] sub_210_d0;
  assign sub_210_d0 = sub_210_s0 - sub_210_s1;
  // sub:221
  wire [16:0] sub_221_s0;
  assign sub_221_s0 = stage_12_pr;
  wire [15:0] sub_221_s1;
  assign sub_221_s1 = di_12;
  wire [16:0] sub_221_d0;
  assign sub_221_d0 = sub_221_s0 - sub_221_s1;
  // sub:232
  wire [16:0] sub_232_s0;
  assign sub_232_s0 = stage_11_pr;
  wire [15:0] sub_232_s1;
  assign sub_232_s1 = di_11;
  wire [16:0] sub_232_d0;
  assign sub_232_d0 = sub_232_s0 - sub_232_s1;
  // sub:243
  wire [16:0] sub_243_s0;
  assign sub_243_s0 = stage_10_pr;
  wire [15:0] sub_243_s1;
  assign sub_243_s1 = di_10;
  wire [16:0] sub_243_d0;
  assign sub_243_d0 = sub_243_s0 - sub_243_s1;
  // sub:254
  wire [16:0] sub_254_s0;
  assign sub_254_s0 = stage_9_pr;
  wire [15:0] sub_254_s1;
  assign sub_254_s1 = di_09;
  wire [16:0] sub_254_d0;
  assign sub_254_d0 = sub_254_s0 - sub_254_s1;
  // sub:265
  wire [16:0] sub_265_s0;
  assign sub_265_s0 = stage_8_pr;
  wire [15:0] sub_265_s1;
  assign sub_265_s1 = di_08;
  wire [16:0] sub_265_d0;
  assign sub_265_d0 = sub_265_s0 - sub_265_s1;
  // sub:276
  wire [16:0] sub_276_s0;
  assign sub_276_s0 = stage_7_pr;
  wire [15:0] sub_276_s1;
  assign sub_276_s1 = di_07;
  wire [16:0] sub_276_d0;
  assign sub_276_d0 = sub_276_s0 - sub_276_s1;
  // sub:287
  wire [16:0] sub_287_s0;
  assign sub_287_s0 = stage_6_pr;
  wire [15:0] sub_287_s1;
  assign sub_287_s1 = di_06;
  wire [16:0] sub_287_d0;
  assign sub_287_d0 = sub_287_s0 - sub_287_s1;
  // sub:298
  wire [16:0] sub_298_s0;
  assign sub_298_s0 = stage_5_pr;
  wire [15:0] sub_298_s1;
  assign sub_298_s1 = di_05;
  wire [16:0] sub_298_d0;
  assign sub_298_d0 = sub_298_s0 - sub_298_s1;
  // sub:309
  wire [16:0] sub_309_s0;
  assign sub_309_s0 = stage_4_pr;
  wire [15:0] sub_309_s1;
  assign sub_309_s1 = di_04;
  wire [16:0] sub_309_d0;
  assign sub_309_d0 = sub_309_s0 - sub_309_s1;
  // sub:320
  wire [16:0] sub_320_s0;
  assign sub_320_s0 = stage_3_pr;
  wire [15:0] sub_320_s1;
  assign sub_320_s1 = di_03;
  wire [16:0] sub_320_d0;
  assign sub_320_d0 = sub_320_s0 - sub_320_s1;
  // sub:331
  wire [16:0] sub_331_s0;
  assign sub_331_s0 = stage_2_pr;
  wire [15:0] sub_331_s1;
  assign sub_331_s1 = di_02;
  wire [16:0] sub_331_d0;
  assign sub_331_d0 = sub_331_s0 - sub_331_s1;
  // sub:342
  wire [16:0] sub_342_s0;
  assign sub_342_s0 = stage_1_pr;
  wire [15:0] sub_342_s1;
  assign sub_342_s1 = di_01;
  wire [16:0] sub_342_d0;
  assign sub_342_d0 = sub_342_s0 - sub_342_s1;
  // sub:353
  wire [16:0] sub_353_s0;
  assign sub_353_s0 = stage_0_pr;
  wire [15:0] sub_353_s1;
  assign sub_353_s1 = di_00;
  wire [16:0] sub_353_d0;
  assign sub_353_d0 = sub_353_s0 - sub_353_s1;
  // Insn wires
  wire  [31:0] insn_o_1_2_0;
  wire  [47:0] insn_o_1_3_0;
  wire  [0:0] insn_o_1_4_0;
  wire  [47:0] insn_o_1_5_0;
  wire  [15:0] insn_o_1_6_0;
  wire  [16:0] insn_o_1_8_0;
  wire  [16:0] insn_o_1_9_0;
  wire  [15:0] insn_o_1_10_0;
  wire  [15:0] insn_o_1_11_0;
  wire  [0:0] insn_o_1_12_0;
  wire  [15:0] insn_o_1_13_0;
  wire  [30:0] insn_o_1_14_0;
  wire  [0:0] insn_o_1_15_0;
  wire  [47:0] insn_o_1_16_0;
  wire  [47:0] insn_o_1_17_0;
  wire  [15:0] insn_o_1_18_0;
  wire  [16:0] insn_o_1_20_0;
  wire  [16:0] insn_o_1_21_0;
  wire  [15:0] insn_o_1_22_0;
  wire  [15:0] insn_o_1_23_0;
  wire  [0:0] insn_o_1_24_0;
  wire  [15:0] insn_o_1_25_0;
  wire  [30:0] insn_o_1_26_0;
  wire  [0:0] insn_o_1_27_0;
  wire  [47:0] insn_o_1_28_0;
  wire  [47:0] insn_o_1_29_0;
  wire  [15:0] insn_o_1_30_0;
  wire  [16:0] insn_o_1_32_0;
  wire  [16:0] insn_o_1_33_0;
  wire  [15:0] insn_o_1_34_0;
  wire  [15:0] insn_o_1_35_0;
  wire  [0:0] insn_o_1_36_0;
  wire  [15:0] insn_o_1_37_0;
  wire  [30:0] insn_o_1_38_0;
  wire  [0:0] insn_o_1_39_0;
  wire  [47:0] insn_o_1_40_0;
  wire  [47:0] insn_o_1_41_0;
  wire  [15:0] insn_o_1_42_0;
  wire  [16:0] insn_o_1_44_0;
  wire  [16:0] insn_o_1_45_0;
  wire  [15:0] insn_o_1_46_0;
  wire  [15:0] insn_o_1_47_0;
  wire  [0:0] insn_o_1_48_0;
  wire  [15:0] insn_o_1_49_0;
  wire  [30:0] insn_o_1_50_0;
  wire  [0:0] insn_o_1_51_0;
  wire  [47:0] insn_o_1_52_0;
  wire  [47:0] insn_o_1_53_0;
  wire  [15:0] insn_o_1_54_0;
  wire  [16:0] insn_o_1_56_0;
  wire  [16:0] insn_o_1_57_0;
  wire  [15:0] insn_o_1_58_0;
  wire  [15:0] insn_o_1_59_0;
  wire  [0:0] insn_o_1_60_0;
  wire  [15:0] insn_o_1_61_0;
  wire  [30:0] insn_o_1_62_0;
  wire  [0:0] insn_o_1_63_0;
  wire  [47:0] insn_o_1_64_0;
  wire  [47:0] insn_o_1_65_0;
  wire  [15:0] insn_o_1_66_0;
  wire  [16:0] insn_o_1_68_0;
  wire  [16:0] insn_o_1_69_0;
  wire  [15:0] insn_o_1_70_0;
  wire  [15:0] insn_o_1_71_0;
  wire  [0:0] insn_o_1_72_0;
  wire  [15:0] insn_o_1_73_0;
  wire  [30:0] insn_o_1_74_0;
  wire  [0:0] insn_o_1_75_0;
  wire  [47:0] insn_o_1_76_0;
  wire  [47:0] insn_o_1_77_0;
  wire  [15:0] insn_o_1_78_0;
  wire  [16:0] insn_o_1_80_0;
  wire  [16:0] insn_o_1_81_0;
  wire  [15:0] insn_o_1_82_0;
  wire  [15:0] insn_o_1_83_0;
  wire  [0:0] insn_o_1_84_0;
  wire  [15:0] insn_o_1_85_0;
  wire  [30:0] insn_o_1_86_0;
  wire  [0:0] insn_o_1_87_0;
  wire  [47:0] insn_o_1_88_0;
  wire  [47:0] insn_o_1_89_0;
  wire  [15:0] insn_o_1_90_0;
  wire  [16:0] insn_o_1_92_0;
  wire  [16:0] insn_o_1_93_0;
  wire  [15:0] insn_o_1_94_0;
  wire  [15:0] insn_o_1_95_0;
  wire  [0:0] insn_o_1_96_0;
  wire  [15:0] insn_o_1_97_0;
  wire  [30:0] insn_o_1_98_0;
  wire  [0:0] insn_o_1_99_0;
  wire  [47:0] insn_o_1_100_0;
  wire  [47:0] insn_o_1_101_0;
  wire  [15:0] insn_o_1_102_0;
  wire  [16:0] insn_o_1_104_0;
  wire  [16:0] insn_o_1_105_0;
  wire  [15:0] insn_o_1_106_0;
  wire  [15:0] insn_o_1_107_0;
  wire  [0:0] insn_o_1_108_0;
  wire  [15:0] insn_o_1_109_0;
  wire  [30:0] insn_o_1_110_0;
  wire  [0:0] insn_o_1_111_0;
  wire  [47:0] insn_o_1_112_0;
  wire  [47:0] insn_o_1_113_0;
  wire  [15:0] insn_o_1_114_0;
  wire  [16:0] insn_o_1_116_0;
  wire  [16:0] insn_o_1_117_0;
  wire  [15:0] insn_o_1_118_0;
  wire  [15:0] insn_o_1_119_0;
  wire  [0:0] insn_o_1_120_0;
  wire  [15:0] insn_o_1_121_0;
  wire  [30:0] insn_o_1_122_0;
  wire  [0:0] insn_o_1_123_0;
  wire  [47:0] insn_o_1_124_0;
  wire  [47:0] insn_o_1_125_0;
  wire  [15:0] insn_o_1_126_0;
  wire  [16:0] insn_o_1_128_0;
  wire  [16:0] insn_o_1_129_0;
  wire  [15:0] insn_o_1_130_0;
  wire  [15:0] insn_o_1_131_0;
  wire  [0:0] insn_o_1_132_0;
  wire  [15:0] insn_o_1_133_0;
  wire  [30:0] insn_o_1_134_0;
  wire  [0:0] insn_o_1_135_0;
  wire  [47:0] insn_o_1_136_0;
  wire  [47:0] insn_o_1_137_0;
  wire  [15:0] insn_o_1_138_0;
  wire  [16:0] insn_o_1_140_0;
  wire  [16:0] insn_o_1_141_0;
  wire  [15:0] insn_o_1_142_0;
  wire  [15:0] insn_o_1_143_0;
  wire  [0:0] insn_o_1_144_0;
  wire  [15:0] insn_o_1_145_0;
  wire  [30:0] insn_o_1_146_0;
  wire  [0:0] insn_o_1_147_0;
  wire  [47:0] insn_o_1_148_0;
  wire  [47:0] insn_o_1_149_0;
  wire  [15:0] insn_o_1_150_0;
  wire  [16:0] insn_o_1_152_0;
  wire  [16:0] insn_o_1_153_0;
  wire  [15:0] insn_o_1_154_0;
  wire  [15:0] insn_o_1_155_0;
  wire  [0:0] insn_o_1_156_0;
  wire  [15:0] insn_o_1_157_0;
  wire  [30:0] insn_o_1_158_0;
  wire  [0:0] insn_o_1_159_0;
  wire  [47:0] insn_o_1_160_0;
  wire  [47:0] insn_o_1_161_0;
  wire  [15:0] insn_o_1_162_0;
  wire  [16:0] insn_o_1_164_0;
  wire  [16:0] insn_o_1_165_0;
  wire  [15:0] insn_o_1_166_0;
  wire  [15:0] insn_o_1_167_0;
  wire  [0:0] insn_o_1_168_0;
  wire  [15:0] insn_o_1_169_0;
  wire  [30:0] insn_o_1_170_0;
  wire  [0:0] insn_o_1_171_0;
  wire  [47:0] insn_o_1_172_0;
  wire  [47:0] insn_o_1_173_0;
  wire  [15:0] insn_o_1_174_0;
  wire  [16:0] insn_o_1_176_0;
  wire  [16:0] insn_o_1_177_0;
  wire  [15:0] insn_o_1_178_0;
  wire  [15:0] insn_o_1_179_0;
  wire  [0:0] insn_o_1_180_0;
  wire  [15:0] insn_o_1_181_0;
  wire  [30:0] insn_o_1_182_0;
  wire  [0:0] insn_o_1_183_0;
  wire  [47:0] insn_o_1_184_0;
  wire  [47:0] insn_o_1_185_0;
  wire  [15:0] insn_o_1_186_0;
  wire  [16:0] insn_o_1_188_0;
  wire  [16:0] insn_o_1_189_0;
  wire  [15:0] insn_o_1_190_0;
  wire  [15:0] insn_o_1_191_0;
  wire  [0:0] insn_o_1_192_0;
  wire  [15:0] insn_o_1_193_0;
  wire  [30:0] insn_o_1_194_0;
  wire  [0:0] insn_o_1_195_0;
  wire  [47:0] insn_o_1_196_0;
  wire  [47:0] insn_o_1_197_0;
  wire  [15:0] insn_o_1_198_0;
  wire  [16:0] insn_o_1_200_0;
  wire  [16:0] insn_o_1_201_0;
  wire  [15:0] insn_o_1_202_0;
  wire  [15:0] insn_o_1_203_0;
  wire  [0:0] insn_o_1_204_0;
  wire  [15:0] insn_o_1_205_0;
  wire  [30:0] insn_o_1_206_0;
  wire  [0:0] insn_o_1_207_0;
  wire  [47:0] insn_o_1_208_0;
  wire  [47:0] insn_o_1_209_0;
  wire  [15:0] insn_o_1_210_0;
  wire  [16:0] insn_o_1_212_0;
  wire  [16:0] insn_o_1_213_0;
  wire  [15:0] insn_o_1_214_0;
  wire  [15:0] insn_o_1_215_0;
  wire  [0:0] insn_o_1_216_0;
  wire  [15:0] insn_o_1_217_0;
  wire  [30:0] insn_o_1_218_0;
  wire  [0:0] insn_o_1_219_0;
  wire  [47:0] insn_o_1_220_0;
  wire  [47:0] insn_o_1_221_0;
  wire  [15:0] insn_o_1_222_0;
  wire  [16:0] insn_o_1_224_0;
  wire  [16:0] insn_o_1_225_0;
  wire  [15:0] insn_o_1_226_0;
  wire  [15:0] insn_o_1_227_0;
  wire  [0:0] insn_o_1_228_0;
  wire  [15:0] insn_o_1_229_0;
  wire  [30:0] insn_o_1_230_0;
  wire  [0:0] insn_o_1_231_0;
  wire  [47:0] insn_o_1_232_0;
  wire  [47:0] insn_o_1_233_0;
  wire  [15:0] insn_o_1_234_0;
  wire  [16:0] insn_o_1_236_0;
  wire  [16:0] insn_o_1_237_0;
  wire  [15:0] insn_o_1_238_0;
  wire  [15:0] insn_o_1_239_0;
  wire  [0:0] insn_o_1_240_0;
  wire  [15:0] insn_o_1_241_0;
  wire  [30:0] insn_o_1_242_0;
  wire  [0:0] insn_o_1_243_0;
  wire  [47:0] insn_o_1_244_0;
  wire  [47:0] insn_o_1_245_0;
  wire  [15:0] insn_o_1_246_0;
  wire  [16:0] insn_o_1_248_0;
  wire  [16:0] insn_o_1_249_0;
  wire  [15:0] insn_o_1_250_0;
  wire  [15:0] insn_o_1_251_0;
  wire  [0:0] insn_o_1_252_0;
  wire  [15:0] insn_o_1_253_0;
  wire  [30:0] insn_o_1_254_0;
  wire  [0:0] insn_o_1_255_0;
  wire  [47:0] insn_o_1_256_0;
  wire  [47:0] insn_o_1_257_0;
  wire  [15:0] insn_o_1_258_0;
  wire  [16:0] insn_o_1_260_0;
  wire  [16:0] insn_o_1_261_0;
  wire  [15:0] insn_o_1_262_0;
  wire  [15:0] insn_o_1_263_0;
  wire  [0:0] insn_o_1_264_0;
  wire  [15:0] insn_o_1_265_0;
  wire  [30:0] insn_o_1_266_0;
  wire  [0:0] insn_o_1_267_0;
  wire  [47:0] insn_o_1_268_0;
  wire  [47:0] insn_o_1_269_0;
  wire  [15:0] insn_o_1_270_0;
  wire  [16:0] insn_o_1_272_0;
  wire  [16:0] insn_o_1_273_0;
  wire  [15:0] insn_o_1_274_0;
  wire  [15:0] insn_o_1_275_0;
  wire  [0:0] insn_o_1_276_0;
  wire  [15:0] insn_o_1_277_0;
  wire  [30:0] insn_o_1_278_0;
  wire  [0:0] insn_o_1_279_0;
  wire  [47:0] insn_o_1_280_0;
  wire  [47:0] insn_o_1_281_0;
  wire  [15:0] insn_o_1_282_0;
  wire  [16:0] insn_o_1_284_0;
  wire  [16:0] insn_o_1_285_0;
  wire  [15:0] insn_o_1_286_0;
  wire  [15:0] insn_o_1_287_0;
  wire  [0:0] insn_o_1_288_0;
  wire  [15:0] insn_o_1_289_0;
  wire  [30:0] insn_o_1_290_0;
  wire  [0:0] insn_o_1_291_0;
  wire  [47:0] insn_o_1_292_0;
  wire  [47:0] insn_o_1_293_0;
  wire  [15:0] insn_o_1_294_0;
  wire  [16:0] insn_o_1_296_0;
  wire  [16:0] insn_o_1_297_0;
  wire  [15:0] insn_o_1_298_0;
  wire  [15:0] insn_o_1_299_0;
  wire  [0:0] insn_o_1_300_0;
  wire  [15:0] insn_o_1_301_0;
  wire  [30:0] insn_o_1_302_0;
  wire  [0:0] insn_o_1_303_0;
  wire  [47:0] insn_o_1_304_0;
  wire  [47:0] insn_o_1_305_0;
  wire  [15:0] insn_o_1_306_0;
  wire  [16:0] insn_o_1_308_0;
  wire  [16:0] insn_o_1_309_0;
  wire  [15:0] insn_o_1_310_0;
  wire  [15:0] insn_o_1_311_0;
  wire  [0:0] insn_o_1_312_0;
  wire  [15:0] insn_o_1_313_0;
  wire  [30:0] insn_o_1_314_0;
  wire  [0:0] insn_o_1_315_0;
  wire  [47:0] insn_o_1_316_0;
  wire  [47:0] insn_o_1_317_0;
  wire  [15:0] insn_o_1_318_0;
  wire  [16:0] insn_o_1_320_0;
  wire  [16:0] insn_o_1_321_0;
  wire  [15:0] insn_o_1_322_0;
  wire  [15:0] insn_o_1_323_0;
  wire  [0:0] insn_o_1_324_0;
  wire  [15:0] insn_o_1_325_0;
  wire  [30:0] insn_o_1_326_0;
  wire  [0:0] insn_o_1_327_0;
  wire  [47:0] insn_o_1_328_0;
  wire  [47:0] insn_o_1_329_0;
  wire  [15:0] insn_o_1_330_0;
  wire  [16:0] insn_o_1_332_0;
  wire  [16:0] insn_o_1_333_0;
  wire  [15:0] insn_o_1_334_0;
  wire  [15:0] insn_o_1_335_0;
  wire  [0:0] insn_o_1_336_0;
  wire  [15:0] insn_o_1_337_0;
  wire  [30:0] insn_o_1_338_0;
  wire  [0:0] insn_o_1_339_0;
  wire  [47:0] insn_o_1_340_0;
  wire  [47:0] insn_o_1_341_0;
  wire  [15:0] insn_o_1_342_0;
  wire  [16:0] insn_o_1_344_0;
  wire  [16:0] insn_o_1_345_0;
  wire  [15:0] insn_o_1_346_0;
  wire  [15:0] insn_o_1_347_0;
  wire  [0:0] insn_o_1_348_0;
  wire  [15:0] insn_o_1_349_0;
  wire  [30:0] insn_o_1_350_0;
  wire  [0:0] insn_o_1_351_0;
  wire  [47:0] insn_o_1_352_0;
  wire  [47:0] insn_o_1_353_0;
  wire  [15:0] insn_o_1_354_0;
  wire  [16:0] insn_o_1_356_0;
  wire  [16:0] insn_o_1_357_0;
  wire  [15:0] insn_o_1_358_0;
  wire  [15:0] insn_o_1_359_0;
  wire  [0:0] insn_o_1_360_0;
  wire  [15:0] insn_o_1_361_0;
  wire  [30:0] insn_o_1_362_0;
  wire  [0:0] insn_o_1_363_0;
  wire  [47:0] insn_o_1_364_0;
  wire  [47:0] insn_o_1_365_0;
  wire  [15:0] insn_o_1_366_0;
  wire  [16:0] insn_o_1_368_0;
  wire  [16:0] insn_o_1_369_0;
  wire  [15:0] insn_o_1_370_0;
  wire  [15:0] insn_o_1_371_0;
  wire  [0:0] insn_o_1_372_0;
  wire  [15:0] insn_o_1_373_0;
  wire  [30:0] insn_o_1_374_0;
  wire  [0:0] insn_o_1_375_0;
  wire  [47:0] insn_o_1_376_0;
  wire  [47:0] insn_o_1_377_0;
  wire  [15:0] insn_o_1_378_0;
  wire  [16:0] insn_o_1_380_0;
  wire  [16:0] insn_o_1_381_0;
  wire  [15:0] insn_o_1_382_0;
  wire  [15:0] insn_o_1_383_0;
  wire  [0:0] insn_o_1_384_0;
  wire  [15:0] insn_o_1_385_0;
  wire  [30:0] insn_o_1_386_0;
  wire  [0:0] insn_o_1_387_0;
  wire  [47:0] insn_o_1_388_0;
  wire  [15:0] insn_o_1_389_0;
  wire  [31:0] insn_o_1_390_0;
  // Insn assigns
  assign insn_o_1_2_0 = dividend;
  assign stage_32_zi_l = insn_o_1_2_0;
  assign insn_o_1_3_0 = {16'd0, stage_32_zi_l};
  assign stage_32_zi_i = insn_o_1_3_0;
  assign insn_o_1_4_0 = i_valid;
  assign start = insn_o_1_4_0;
  assign insn_o_1_6_0 = divisor;
  assign insn_o_1_8_0 = zi_31[47:31];
  assign stage_31_pr = insn_o_1_8_0;
  assign insn_o_1_9_0 = sub_12_d0;
  assign stage_31_sb = insn_o_1_9_0;
  assign insn_o_1_10_0 = stage_31_sb[15:0];
  assign stage_31_m0 = insn_o_1_10_0;
  assign insn_o_1_11_0 = stage_31_pr[15:0];
  assign stage_31_m1 = insn_o_1_11_0;
  assign insn_o_1_12_0 = stage_31_sb[16:16];
  assign stage_31_ms = insn_o_1_12_0;
  assign insn_o_1_13_0 = stage_31_ms ? stage_31_m1 : stage_31_m0;
  assign stage_31_mx = insn_o_1_13_0;
  assign insn_o_1_14_0 = zi_31[30:0];
  assign stage_31_zl = insn_o_1_14_0;
  assign insn_o_1_15_0 = ~stage_31_ms;
  assign stage_31_zb = insn_o_1_15_0;
  assign insn_o_1_16_0 = {stage_31_mx, stage_31_zl, stage_31_zb};
  assign stage_31_zo = insn_o_1_16_0;
  assign insn_o_1_20_0 = zi_30[47:31];
  assign stage_30_pr = insn_o_1_20_0;
  assign insn_o_1_21_0 = sub_23_d0;
  assign stage_30_sb = insn_o_1_21_0;
  assign insn_o_1_22_0 = stage_30_sb[15:0];
  assign stage_30_m0 = insn_o_1_22_0;
  assign insn_o_1_23_0 = stage_30_pr[15:0];
  assign stage_30_m1 = insn_o_1_23_0;
  assign insn_o_1_24_0 = stage_30_sb[16:16];
  assign stage_30_ms = insn_o_1_24_0;
  assign insn_o_1_25_0 = stage_30_ms ? stage_30_m1 : stage_30_m0;
  assign stage_30_mx = insn_o_1_25_0;
  assign insn_o_1_26_0 = zi_30[30:0];
  assign stage_30_zl = insn_o_1_26_0;
  assign insn_o_1_27_0 = ~stage_30_ms;
  assign stage_30_zb = insn_o_1_27_0;
  assign insn_o_1_28_0 = {stage_30_mx, stage_30_zl, stage_30_zb};
  assign stage_30_zo = insn_o_1_28_0;
  assign insn_o_1_32_0 = zi_29[47:31];
  assign stage_29_pr = insn_o_1_32_0;
  assign insn_o_1_33_0 = sub_34_d0;
  assign stage_29_sb = insn_o_1_33_0;
  assign insn_o_1_34_0 = stage_29_sb[15:0];
  assign stage_29_m0 = insn_o_1_34_0;
  assign insn_o_1_35_0 = stage_29_pr[15:0];
  assign stage_29_m1 = insn_o_1_35_0;
  assign insn_o_1_36_0 = stage_29_sb[16:16];
  assign stage_29_ms = insn_o_1_36_0;
  assign insn_o_1_37_0 = stage_29_ms ? stage_29_m1 : stage_29_m0;
  assign stage_29_mx = insn_o_1_37_0;
  assign insn_o_1_38_0 = zi_29[30:0];
  assign stage_29_zl = insn_o_1_38_0;
  assign insn_o_1_39_0 = ~stage_29_ms;
  assign stage_29_zb = insn_o_1_39_0;
  assign insn_o_1_40_0 = {stage_29_mx, stage_29_zl, stage_29_zb};
  assign stage_29_zo = insn_o_1_40_0;
  assign insn_o_1_44_0 = zi_28[47:31];
  assign stage_28_pr = insn_o_1_44_0;
  assign insn_o_1_45_0 = sub_45_d0;
  assign stage_28_sb = insn_o_1_45_0;
  assign insn_o_1_46_0 = stage_28_sb[15:0];
  assign stage_28_m0 = insn_o_1_46_0;
  assign insn_o_1_47_0 = stage_28_pr[15:0];
  assign stage_28_m1 = insn_o_1_47_0;
  assign insn_o_1_48_0 = stage_28_sb[16:16];
  assign stage_28_ms = insn_o_1_48_0;
  assign insn_o_1_49_0 = stage_28_ms ? stage_28_m1 : stage_28_m0;
  assign stage_28_mx = insn_o_1_49_0;
  assign insn_o_1_50_0 = zi_28[30:0];
  assign stage_28_zl = insn_o_1_50_0;
  assign insn_o_1_51_0 = ~stage_28_ms;
  assign stage_28_zb = insn_o_1_51_0;
  assign insn_o_1_52_0 = {stage_28_mx, stage_28_zl, stage_28_zb};
  assign stage_28_zo = insn_o_1_52_0;
  assign insn_o_1_56_0 = zi_27[47:31];
  assign stage_27_pr = insn_o_1_56_0;
  assign insn_o_1_57_0 = sub_56_d0;
  assign stage_27_sb = insn_o_1_57_0;
  assign insn_o_1_58_0 = stage_27_sb[15:0];
  assign stage_27_m0 = insn_o_1_58_0;
  assign insn_o_1_59_0 = stage_27_pr[15:0];
  assign stage_27_m1 = insn_o_1_59_0;
  assign insn_o_1_60_0 = stage_27_sb[16:16];
  assign stage_27_ms = insn_o_1_60_0;
  assign insn_o_1_61_0 = stage_27_ms ? stage_27_m1 : stage_27_m0;
  assign stage_27_mx = insn_o_1_61_0;
  assign insn_o_1_62_0 = zi_27[30:0];
  assign stage_27_zl = insn_o_1_62_0;
  assign insn_o_1_63_0 = ~stage_27_ms;
  assign stage_27_zb = insn_o_1_63_0;
  assign insn_o_1_64_0 = {stage_27_mx, stage_27_zl, stage_27_zb};
  assign stage_27_zo = insn_o_1_64_0;
  assign insn_o_1_68_0 = zi_26[47:31];
  assign stage_26_pr = insn_o_1_68_0;
  assign insn_o_1_69_0 = sub_67_d0;
  assign stage_26_sb = insn_o_1_69_0;
  assign insn_o_1_70_0 = stage_26_sb[15:0];
  assign stage_26_m0 = insn_o_1_70_0;
  assign insn_o_1_71_0 = stage_26_pr[15:0];
  assign stage_26_m1 = insn_o_1_71_0;
  assign insn_o_1_72_0 = stage_26_sb[16:16];
  assign stage_26_ms = insn_o_1_72_0;
  assign insn_o_1_73_0 = stage_26_ms ? stage_26_m1 : stage_26_m0;
  assign stage_26_mx = insn_o_1_73_0;
  assign insn_o_1_74_0 = zi_26[30:0];
  assign stage_26_zl = insn_o_1_74_0;
  assign insn_o_1_75_0 = ~stage_26_ms;
  assign stage_26_zb = insn_o_1_75_0;
  assign insn_o_1_76_0 = {stage_26_mx, stage_26_zl, stage_26_zb};
  assign stage_26_zo = insn_o_1_76_0;
  assign insn_o_1_80_0 = zi_25[47:31];
  assign stage_25_pr = insn_o_1_80_0;
  assign insn_o_1_81_0 = sub_78_d0;
  assign stage_25_sb = insn_o_1_81_0;
  assign insn_o_1_82_0 = stage_25_sb[15:0];
  assign stage_25_m0 = insn_o_1_82_0;
  assign insn_o_1_83_0 = stage_25_pr[15:0];
  assign stage_25_m1 = insn_o_1_83_0;
  assign insn_o_1_84_0 = stage_25_sb[16:16];
  assign stage_25_ms = insn_o_1_84_0;
  assign insn_o_1_85_0 = stage_25_ms ? stage_25_m1 : stage_25_m0;
  assign stage_25_mx = insn_o_1_85_0;
  assign insn_o_1_86_0 = zi_25[30:0];
  assign stage_25_zl = insn_o_1_86_0;
  assign insn_o_1_87_0 = ~stage_25_ms;
  assign stage_25_zb = insn_o_1_87_0;
  assign insn_o_1_88_0 = {stage_25_mx, stage_25_zl, stage_25_zb};
  assign stage_25_zo = insn_o_1_88_0;
  assign insn_o_1_92_0 = zi_24[47:31];
  assign stage_24_pr = insn_o_1_92_0;
  assign insn_o_1_93_0 = sub_89_d0;
  assign stage_24_sb = insn_o_1_93_0;
  assign insn_o_1_94_0 = stage_24_sb[15:0];
  assign stage_24_m0 = insn_o_1_94_0;
  assign insn_o_1_95_0 = stage_24_pr[15:0];
  assign stage_24_m1 = insn_o_1_95_0;
  assign insn_o_1_96_0 = stage_24_sb[16:16];
  assign stage_24_ms = insn_o_1_96_0;
  assign insn_o_1_97_0 = stage_24_ms ? stage_24_m1 : stage_24_m0;
  assign stage_24_mx = insn_o_1_97_0;
  assign insn_o_1_98_0 = zi_24[30:0];
  assign stage_24_zl = insn_o_1_98_0;
  assign insn_o_1_99_0 = ~stage_24_ms;
  assign stage_24_zb = insn_o_1_99_0;
  assign insn_o_1_100_0 = {stage_24_mx, stage_24_zl, stage_24_zb};
  assign stage_24_zo = insn_o_1_100_0;
  assign insn_o_1_104_0 = zi_23[47:31];
  assign stage_23_pr = insn_o_1_104_0;
  assign insn_o_1_105_0 = sub_100_d0;
  assign stage_23_sb = insn_o_1_105_0;
  assign insn_o_1_106_0 = stage_23_sb[15:0];
  assign stage_23_m0 = insn_o_1_106_0;
  assign insn_o_1_107_0 = stage_23_pr[15:0];
  assign stage_23_m1 = insn_o_1_107_0;
  assign insn_o_1_108_0 = stage_23_sb[16:16];
  assign stage_23_ms = insn_o_1_108_0;
  assign insn_o_1_109_0 = stage_23_ms ? stage_23_m1 : stage_23_m0;
  assign stage_23_mx = insn_o_1_109_0;
  assign insn_o_1_110_0 = zi_23[30:0];
  assign stage_23_zl = insn_o_1_110_0;
  assign insn_o_1_111_0 = ~stage_23_ms;
  assign stage_23_zb = insn_o_1_111_0;
  assign insn_o_1_112_0 = {stage_23_mx, stage_23_zl, stage_23_zb};
  assign stage_23_zo = insn_o_1_112_0;
  assign insn_o_1_116_0 = zi_22[47:31];
  assign stage_22_pr = insn_o_1_116_0;
  assign insn_o_1_117_0 = sub_111_d0;
  assign stage_22_sb = insn_o_1_117_0;
  assign insn_o_1_118_0 = stage_22_sb[15:0];
  assign stage_22_m0 = insn_o_1_118_0;
  assign insn_o_1_119_0 = stage_22_pr[15:0];
  assign stage_22_m1 = insn_o_1_119_0;
  assign insn_o_1_120_0 = stage_22_sb[16:16];
  assign stage_22_ms = insn_o_1_120_0;
  assign insn_o_1_121_0 = stage_22_ms ? stage_22_m1 : stage_22_m0;
  assign stage_22_mx = insn_o_1_121_0;
  assign insn_o_1_122_0 = zi_22[30:0];
  assign stage_22_zl = insn_o_1_122_0;
  assign insn_o_1_123_0 = ~stage_22_ms;
  assign stage_22_zb = insn_o_1_123_0;
  assign insn_o_1_124_0 = {stage_22_mx, stage_22_zl, stage_22_zb};
  assign stage_22_zo = insn_o_1_124_0;
  assign insn_o_1_128_0 = zi_21[47:31];
  assign stage_21_pr = insn_o_1_128_0;
  assign insn_o_1_129_0 = sub_122_d0;
  assign stage_21_sb = insn_o_1_129_0;
  assign insn_o_1_130_0 = stage_21_sb[15:0];
  assign stage_21_m0 = insn_o_1_130_0;
  assign insn_o_1_131_0 = stage_21_pr[15:0];
  assign stage_21_m1 = insn_o_1_131_0;
  assign insn_o_1_132_0 = stage_21_sb[16:16];
  assign stage_21_ms = insn_o_1_132_0;
  assign insn_o_1_133_0 = stage_21_ms ? stage_21_m1 : stage_21_m0;
  assign stage_21_mx = insn_o_1_133_0;
  assign insn_o_1_134_0 = zi_21[30:0];
  assign stage_21_zl = insn_o_1_134_0;
  assign insn_o_1_135_0 = ~stage_21_ms;
  assign stage_21_zb = insn_o_1_135_0;
  assign insn_o_1_136_0 = {stage_21_mx, stage_21_zl, stage_21_zb};
  assign stage_21_zo = insn_o_1_136_0;
  assign insn_o_1_140_0 = zi_20[47:31];
  assign stage_20_pr = insn_o_1_140_0;
  assign insn_o_1_141_0 = sub_133_d0;
  assign stage_20_sb = insn_o_1_141_0;
  assign insn_o_1_142_0 = stage_20_sb[15:0];
  assign stage_20_m0 = insn_o_1_142_0;
  assign insn_o_1_143_0 = stage_20_pr[15:0];
  assign stage_20_m1 = insn_o_1_143_0;
  assign insn_o_1_144_0 = stage_20_sb[16:16];
  assign stage_20_ms = insn_o_1_144_0;
  assign insn_o_1_145_0 = stage_20_ms ? stage_20_m1 : stage_20_m0;
  assign stage_20_mx = insn_o_1_145_0;
  assign insn_o_1_146_0 = zi_20[30:0];
  assign stage_20_zl = insn_o_1_146_0;
  assign insn_o_1_147_0 = ~stage_20_ms;
  assign stage_20_zb = insn_o_1_147_0;
  assign insn_o_1_148_0 = {stage_20_mx, stage_20_zl, stage_20_zb};
  assign stage_20_zo = insn_o_1_148_0;
  assign insn_o_1_152_0 = zi_19[47:31];
  assign stage_19_pr = insn_o_1_152_0;
  assign insn_o_1_153_0 = sub_144_d0;
  assign stage_19_sb = insn_o_1_153_0;
  assign insn_o_1_154_0 = stage_19_sb[15:0];
  assign stage_19_m0 = insn_o_1_154_0;
  assign insn_o_1_155_0 = stage_19_pr[15:0];
  assign stage_19_m1 = insn_o_1_155_0;
  assign insn_o_1_156_0 = stage_19_sb[16:16];
  assign stage_19_ms = insn_o_1_156_0;
  assign insn_o_1_157_0 = stage_19_ms ? stage_19_m1 : stage_19_m0;
  assign stage_19_mx = insn_o_1_157_0;
  assign insn_o_1_158_0 = zi_19[30:0];
  assign stage_19_zl = insn_o_1_158_0;
  assign insn_o_1_159_0 = ~stage_19_ms;
  assign stage_19_zb = insn_o_1_159_0;
  assign insn_o_1_160_0 = {stage_19_mx, stage_19_zl, stage_19_zb};
  assign stage_19_zo = insn_o_1_160_0;
  assign insn_o_1_164_0 = zi_18[47:31];
  assign stage_18_pr = insn_o_1_164_0;
  assign insn_o_1_165_0 = sub_155_d0;
  assign stage_18_sb = insn_o_1_165_0;
  assign insn_o_1_166_0 = stage_18_sb[15:0];
  assign stage_18_m0 = insn_o_1_166_0;
  assign insn_o_1_167_0 = stage_18_pr[15:0];
  assign stage_18_m1 = insn_o_1_167_0;
  assign insn_o_1_168_0 = stage_18_sb[16:16];
  assign stage_18_ms = insn_o_1_168_0;
  assign insn_o_1_169_0 = stage_18_ms ? stage_18_m1 : stage_18_m0;
  assign stage_18_mx = insn_o_1_169_0;
  assign insn_o_1_170_0 = zi_18[30:0];
  assign stage_18_zl = insn_o_1_170_0;
  assign insn_o_1_171_0 = ~stage_18_ms;
  assign stage_18_zb = insn_o_1_171_0;
  assign insn_o_1_172_0 = {stage_18_mx, stage_18_zl, stage_18_zb};
  assign stage_18_zo = insn_o_1_172_0;
  assign insn_o_1_176_0 = zi_17[47:31];
  assign stage_17_pr = insn_o_1_176_0;
  assign insn_o_1_177_0 = sub_166_d0;
  assign stage_17_sb = insn_o_1_177_0;
  assign insn_o_1_178_0 = stage_17_sb[15:0];
  assign stage_17_m0 = insn_o_1_178_0;
  assign insn_o_1_179_0 = stage_17_pr[15:0];
  assign stage_17_m1 = insn_o_1_179_0;
  assign insn_o_1_180_0 = stage_17_sb[16:16];
  assign stage_17_ms = insn_o_1_180_0;
  assign insn_o_1_181_0 = stage_17_ms ? stage_17_m1 : stage_17_m0;
  assign stage_17_mx = insn_o_1_181_0;
  assign insn_o_1_182_0 = zi_17[30:0];
  assign stage_17_zl = insn_o_1_182_0;
  assign insn_o_1_183_0 = ~stage_17_ms;
  assign stage_17_zb = insn_o_1_183_0;
  assign insn_o_1_184_0 = {stage_17_mx, stage_17_zl, stage_17_zb};
  assign stage_17_zo = insn_o_1_184_0;
  assign insn_o_1_188_0 = zi_16[47:31];
  assign stage_16_pr = insn_o_1_188_0;
  assign insn_o_1_189_0 = sub_177_d0;
  assign stage_16_sb = insn_o_1_189_0;
  assign insn_o_1_190_0 = stage_16_sb[15:0];
  assign stage_16_m0 = insn_o_1_190_0;
  assign insn_o_1_191_0 = stage_16_pr[15:0];
  assign stage_16_m1 = insn_o_1_191_0;
  assign insn_o_1_192_0 = stage_16_sb[16:16];
  assign stage_16_ms = insn_o_1_192_0;
  assign insn_o_1_193_0 = stage_16_ms ? stage_16_m1 : stage_16_m0;
  assign stage_16_mx = insn_o_1_193_0;
  assign insn_o_1_194_0 = zi_16[30:0];
  assign stage_16_zl = insn_o_1_194_0;
  assign insn_o_1_195_0 = ~stage_16_ms;
  assign stage_16_zb = insn_o_1_195_0;
  assign insn_o_1_196_0 = {stage_16_mx, stage_16_zl, stage_16_zb};
  assign stage_16_zo = insn_o_1_196_0;
  assign insn_o_1_200_0 = zi_15[47:31];
  assign stage_15_pr = insn_o_1_200_0;
  assign insn_o_1_201_0 = sub_188_d0;
  assign stage_15_sb = insn_o_1_201_0;
  assign insn_o_1_202_0 = stage_15_sb[15:0];
  assign stage_15_m0 = insn_o_1_202_0;
  assign insn_o_1_203_0 = stage_15_pr[15:0];
  assign stage_15_m1 = insn_o_1_203_0;
  assign insn_o_1_204_0 = stage_15_sb[16:16];
  assign stage_15_ms = insn_o_1_204_0;
  assign insn_o_1_205_0 = stage_15_ms ? stage_15_m1 : stage_15_m0;
  assign stage_15_mx = insn_o_1_205_0;
  assign insn_o_1_206_0 = zi_15[30:0];
  assign stage_15_zl = insn_o_1_206_0;
  assign insn_o_1_207_0 = ~stage_15_ms;
  assign stage_15_zb = insn_o_1_207_0;
  assign insn_o_1_208_0 = {stage_15_mx, stage_15_zl, stage_15_zb};
  assign stage_15_zo = insn_o_1_208_0;
  assign insn_o_1_212_0 = zi_14[47:31];
  assign stage_14_pr = insn_o_1_212_0;
  assign insn_o_1_213_0 = sub_199_d0;
  assign stage_14_sb = insn_o_1_213_0;
  assign insn_o_1_214_0 = stage_14_sb[15:0];
  assign stage_14_m0 = insn_o_1_214_0;
  assign insn_o_1_215_0 = stage_14_pr[15:0];
  assign stage_14_m1 = insn_o_1_215_0;
  assign insn_o_1_216_0 = stage_14_sb[16:16];
  assign stage_14_ms = insn_o_1_216_0;
  assign insn_o_1_217_0 = stage_14_ms ? stage_14_m1 : stage_14_m0;
  assign stage_14_mx = insn_o_1_217_0;
  assign insn_o_1_218_0 = zi_14[30:0];
  assign stage_14_zl = insn_o_1_218_0;
  assign insn_o_1_219_0 = ~stage_14_ms;
  assign stage_14_zb = insn_o_1_219_0;
  assign insn_o_1_220_0 = {stage_14_mx, stage_14_zl, stage_14_zb};
  assign stage_14_zo = insn_o_1_220_0;
  assign insn_o_1_224_0 = zi_13[47:31];
  assign stage_13_pr = insn_o_1_224_0;
  assign insn_o_1_225_0 = sub_210_d0;
  assign stage_13_sb = insn_o_1_225_0;
  assign insn_o_1_226_0 = stage_13_sb[15:0];
  assign stage_13_m0 = insn_o_1_226_0;
  assign insn_o_1_227_0 = stage_13_pr[15:0];
  assign stage_13_m1 = insn_o_1_227_0;
  assign insn_o_1_228_0 = stage_13_sb[16:16];
  assign stage_13_ms = insn_o_1_228_0;
  assign insn_o_1_229_0 = stage_13_ms ? stage_13_m1 : stage_13_m0;
  assign stage_13_mx = insn_o_1_229_0;
  assign insn_o_1_230_0 = zi_13[30:0];
  assign stage_13_zl = insn_o_1_230_0;
  assign insn_o_1_231_0 = ~stage_13_ms;
  assign stage_13_zb = insn_o_1_231_0;
  assign insn_o_1_232_0 = {stage_13_mx, stage_13_zl, stage_13_zb};
  assign stage_13_zo = insn_o_1_232_0;
  assign insn_o_1_236_0 = zi_12[47:31];
  assign stage_12_pr = insn_o_1_236_0;
  assign insn_o_1_237_0 = sub_221_d0;
  assign stage_12_sb = insn_o_1_237_0;
  assign insn_o_1_238_0 = stage_12_sb[15:0];
  assign stage_12_m0 = insn_o_1_238_0;
  assign insn_o_1_239_0 = stage_12_pr[15:0];
  assign stage_12_m1 = insn_o_1_239_0;
  assign insn_o_1_240_0 = stage_12_sb[16:16];
  assign stage_12_ms = insn_o_1_240_0;
  assign insn_o_1_241_0 = stage_12_ms ? stage_12_m1 : stage_12_m0;
  assign stage_12_mx = insn_o_1_241_0;
  assign insn_o_1_242_0 = zi_12[30:0];
  assign stage_12_zl = insn_o_1_242_0;
  assign insn_o_1_243_0 = ~stage_12_ms;
  assign stage_12_zb = insn_o_1_243_0;
  assign insn_o_1_244_0 = {stage_12_mx, stage_12_zl, stage_12_zb};
  assign stage_12_zo = insn_o_1_244_0;
  assign insn_o_1_248_0 = zi_11[47:31];
  assign stage_11_pr = insn_o_1_248_0;
  assign insn_o_1_249_0 = sub_232_d0;
  assign stage_11_sb = insn_o_1_249_0;
  assign insn_o_1_250_0 = stage_11_sb[15:0];
  assign stage_11_m0 = insn_o_1_250_0;
  assign insn_o_1_251_0 = stage_11_pr[15:0];
  assign stage_11_m1 = insn_o_1_251_0;
  assign insn_o_1_252_0 = stage_11_sb[16:16];
  assign stage_11_ms = insn_o_1_252_0;
  assign insn_o_1_253_0 = stage_11_ms ? stage_11_m1 : stage_11_m0;
  assign stage_11_mx = insn_o_1_253_0;
  assign insn_o_1_254_0 = zi_11[30:0];
  assign stage_11_zl = insn_o_1_254_0;
  assign insn_o_1_255_0 = ~stage_11_ms;
  assign stage_11_zb = insn_o_1_255_0;
  assign insn_o_1_256_0 = {stage_11_mx, stage_11_zl, stage_11_zb};
  assign stage_11_zo = insn_o_1_256_0;
  assign insn_o_1_260_0 = zi_10[47:31];
  assign stage_10_pr = insn_o_1_260_0;
  assign insn_o_1_261_0 = sub_243_d0;
  assign stage_10_sb = insn_o_1_261_0;
  assign insn_o_1_262_0 = stage_10_sb[15:0];
  assign stage_10_m0 = insn_o_1_262_0;
  assign insn_o_1_263_0 = stage_10_pr[15:0];
  assign stage_10_m1 = insn_o_1_263_0;
  assign insn_o_1_264_0 = stage_10_sb[16:16];
  assign stage_10_ms = insn_o_1_264_0;
  assign insn_o_1_265_0 = stage_10_ms ? stage_10_m1 : stage_10_m0;
  assign stage_10_mx = insn_o_1_265_0;
  assign insn_o_1_266_0 = zi_10[30:0];
  assign stage_10_zl = insn_o_1_266_0;
  assign insn_o_1_267_0 = ~stage_10_ms;
  assign stage_10_zb = insn_o_1_267_0;
  assign insn_o_1_268_0 = {stage_10_mx, stage_10_zl, stage_10_zb};
  assign stage_10_zo = insn_o_1_268_0;
  assign insn_o_1_272_0 = zi_09[47:31];
  assign stage_9_pr = insn_o_1_272_0;
  assign insn_o_1_273_0 = sub_254_d0;
  assign stage_9_sb = insn_o_1_273_0;
  assign insn_o_1_274_0 = stage_9_sb[15:0];
  assign stage_9_m0 = insn_o_1_274_0;
  assign insn_o_1_275_0 = stage_9_pr[15:0];
  assign stage_9_m1 = insn_o_1_275_0;
  assign insn_o_1_276_0 = stage_9_sb[16:16];
  assign stage_9_ms = insn_o_1_276_0;
  assign insn_o_1_277_0 = stage_9_ms ? stage_9_m1 : stage_9_m0;
  assign stage_9_mx = insn_o_1_277_0;
  assign insn_o_1_278_0 = zi_09[30:0];
  assign stage_9_zl = insn_o_1_278_0;
  assign insn_o_1_279_0 = ~stage_9_ms;
  assign stage_9_zb = insn_o_1_279_0;
  assign insn_o_1_280_0 = {stage_9_mx, stage_9_zl, stage_9_zb};
  assign stage_9_zo = insn_o_1_280_0;
  assign insn_o_1_284_0 = zi_08[47:31];
  assign stage_8_pr = insn_o_1_284_0;
  assign insn_o_1_285_0 = sub_265_d0;
  assign stage_8_sb = insn_o_1_285_0;
  assign insn_o_1_286_0 = stage_8_sb[15:0];
  assign stage_8_m0 = insn_o_1_286_0;
  assign insn_o_1_287_0 = stage_8_pr[15:0];
  assign stage_8_m1 = insn_o_1_287_0;
  assign insn_o_1_288_0 = stage_8_sb[16:16];
  assign stage_8_ms = insn_o_1_288_0;
  assign insn_o_1_289_0 = stage_8_ms ? stage_8_m1 : stage_8_m0;
  assign stage_8_mx = insn_o_1_289_0;
  assign insn_o_1_290_0 = zi_08[30:0];
  assign stage_8_zl = insn_o_1_290_0;
  assign insn_o_1_291_0 = ~stage_8_ms;
  assign stage_8_zb = insn_o_1_291_0;
  assign insn_o_1_292_0 = {stage_8_mx, stage_8_zl, stage_8_zb};
  assign stage_8_zo = insn_o_1_292_0;
  assign insn_o_1_296_0 = zi_07[47:31];
  assign stage_7_pr = insn_o_1_296_0;
  assign insn_o_1_297_0 = sub_276_d0;
  assign stage_7_sb = insn_o_1_297_0;
  assign insn_o_1_298_0 = stage_7_sb[15:0];
  assign stage_7_m0 = insn_o_1_298_0;
  assign insn_o_1_299_0 = stage_7_pr[15:0];
  assign stage_7_m1 = insn_o_1_299_0;
  assign insn_o_1_300_0 = stage_7_sb[16:16];
  assign stage_7_ms = insn_o_1_300_0;
  assign insn_o_1_301_0 = stage_7_ms ? stage_7_m1 : stage_7_m0;
  assign stage_7_mx = insn_o_1_301_0;
  assign insn_o_1_302_0 = zi_07[30:0];
  assign stage_7_zl = insn_o_1_302_0;
  assign insn_o_1_303_0 = ~stage_7_ms;
  assign stage_7_zb = insn_o_1_303_0;
  assign insn_o_1_304_0 = {stage_7_mx, stage_7_zl, stage_7_zb};
  assign stage_7_zo = insn_o_1_304_0;
  assign insn_o_1_308_0 = zi_06[47:31];
  assign stage_6_pr = insn_o_1_308_0;
  assign insn_o_1_309_0 = sub_287_d0;
  assign stage_6_sb = insn_o_1_309_0;
  assign insn_o_1_310_0 = stage_6_sb[15:0];
  assign stage_6_m0 = insn_o_1_310_0;
  assign insn_o_1_311_0 = stage_6_pr[15:0];
  assign stage_6_m1 = insn_o_1_311_0;
  assign insn_o_1_312_0 = stage_6_sb[16:16];
  assign stage_6_ms = insn_o_1_312_0;
  assign insn_o_1_313_0 = stage_6_ms ? stage_6_m1 : stage_6_m0;
  assign stage_6_mx = insn_o_1_313_0;
  assign insn_o_1_314_0 = zi_06[30:0];
  assign stage_6_zl = insn_o_1_314_0;
  assign insn_o_1_315_0 = ~stage_6_ms;
  assign stage_6_zb = insn_o_1_315_0;
  assign insn_o_1_316_0 = {stage_6_mx, stage_6_zl, stage_6_zb};
  assign stage_6_zo = insn_o_1_316_0;
  assign insn_o_1_320_0 = zi_05[47:31];
  assign stage_5_pr = insn_o_1_320_0;
  assign insn_o_1_321_0 = sub_298_d0;
  assign stage_5_sb = insn_o_1_321_0;
  assign insn_o_1_322_0 = stage_5_sb[15:0];
  assign stage_5_m0 = insn_o_1_322_0;
  assign insn_o_1_323_0 = stage_5_pr[15:0];
  assign stage_5_m1 = insn_o_1_323_0;
  assign insn_o_1_324_0 = stage_5_sb[16:16];
  assign stage_5_ms = insn_o_1_324_0;
  assign insn_o_1_325_0 = stage_5_ms ? stage_5_m1 : stage_5_m0;
  assign stage_5_mx = insn_o_1_325_0;
  assign insn_o_1_326_0 = zi_05[30:0];
  assign stage_5_zl = insn_o_1_326_0;
  assign insn_o_1_327_0 = ~stage_5_ms;
  assign stage_5_zb = insn_o_1_327_0;
  assign insn_o_1_328_0 = {stage_5_mx, stage_5_zl, stage_5_zb};
  assign stage_5_zo = insn_o_1_328_0;
  assign insn_o_1_332_0 = zi_04[47:31];
  assign stage_4_pr = insn_o_1_332_0;
  assign insn_o_1_333_0 = sub_309_d0;
  assign stage_4_sb = insn_o_1_333_0;
  assign insn_o_1_334_0 = stage_4_sb[15:0];
  assign stage_4_m0 = insn_o_1_334_0;
  assign insn_o_1_335_0 = stage_4_pr[15:0];
  assign stage_4_m1 = insn_o_1_335_0;
  assign insn_o_1_336_0 = stage_4_sb[16:16];
  assign stage_4_ms = insn_o_1_336_0;
  assign insn_o_1_337_0 = stage_4_ms ? stage_4_m1 : stage_4_m0;
  assign stage_4_mx = insn_o_1_337_0;
  assign insn_o_1_338_0 = zi_04[30:0];
  assign stage_4_zl = insn_o_1_338_0;
  assign insn_o_1_339_0 = ~stage_4_ms;
  assign stage_4_zb = insn_o_1_339_0;
  assign insn_o_1_340_0 = {stage_4_mx, stage_4_zl, stage_4_zb};
  assign stage_4_zo = insn_o_1_340_0;
  assign insn_o_1_344_0 = zi_03[47:31];
  assign stage_3_pr = insn_o_1_344_0;
  assign insn_o_1_345_0 = sub_320_d0;
  assign stage_3_sb = insn_o_1_345_0;
  assign insn_o_1_346_0 = stage_3_sb[15:0];
  assign stage_3_m0 = insn_o_1_346_0;
  assign insn_o_1_347_0 = stage_3_pr[15:0];
  assign stage_3_m1 = insn_o_1_347_0;
  assign insn_o_1_348_0 = stage_3_sb[16:16];
  assign stage_3_ms = insn_o_1_348_0;
  assign insn_o_1_349_0 = stage_3_ms ? stage_3_m1 : stage_3_m0;
  assign stage_3_mx = insn_o_1_349_0;
  assign insn_o_1_350_0 = zi_03[30:0];
  assign stage_3_zl = insn_o_1_350_0;
  assign insn_o_1_351_0 = ~stage_3_ms;
  assign stage_3_zb = insn_o_1_351_0;
  assign insn_o_1_352_0 = {stage_3_mx, stage_3_zl, stage_3_zb};
  assign stage_3_zo = insn_o_1_352_0;
  assign insn_o_1_356_0 = zi_02[47:31];
  assign stage_2_pr = insn_o_1_356_0;
  assign insn_o_1_357_0 = sub_331_d0;
  assign stage_2_sb = insn_o_1_357_0;
  assign insn_o_1_358_0 = stage_2_sb[15:0];
  assign stage_2_m0 = insn_o_1_358_0;
  assign insn_o_1_359_0 = stage_2_pr[15:0];
  assign stage_2_m1 = insn_o_1_359_0;
  assign insn_o_1_360_0 = stage_2_sb[16:16];
  assign stage_2_ms = insn_o_1_360_0;
  assign insn_o_1_361_0 = stage_2_ms ? stage_2_m1 : stage_2_m0;
  assign stage_2_mx = insn_o_1_361_0;
  assign insn_o_1_362_0 = zi_02[30:0];
  assign stage_2_zl = insn_o_1_362_0;
  assign insn_o_1_363_0 = ~stage_2_ms;
  assign stage_2_zb = insn_o_1_363_0;
  assign insn_o_1_364_0 = {stage_2_mx, stage_2_zl, stage_2_zb};
  assign stage_2_zo = insn_o_1_364_0;
  assign insn_o_1_368_0 = zi_01[47:31];
  assign stage_1_pr = insn_o_1_368_0;
  assign insn_o_1_369_0 = sub_342_d0;
  assign stage_1_sb = insn_o_1_369_0;
  assign insn_o_1_370_0 = stage_1_sb[15:0];
  assign stage_1_m0 = insn_o_1_370_0;
  assign insn_o_1_371_0 = stage_1_pr[15:0];
  assign stage_1_m1 = insn_o_1_371_0;
  assign insn_o_1_372_0 = stage_1_sb[16:16];
  assign stage_1_ms = insn_o_1_372_0;
  assign insn_o_1_373_0 = stage_1_ms ? stage_1_m1 : stage_1_m0;
  assign stage_1_mx = insn_o_1_373_0;
  assign insn_o_1_374_0 = zi_01[30:0];
  assign stage_1_zl = insn_o_1_374_0;
  assign insn_o_1_375_0 = ~stage_1_ms;
  assign stage_1_zb = insn_o_1_375_0;
  assign insn_o_1_376_0 = {stage_1_mx, stage_1_zl, stage_1_zb};
  assign stage_1_zo = insn_o_1_376_0;
  assign insn_o_1_380_0 = zi_00[47:31];
  assign stage_0_pr = insn_o_1_380_0;
  assign insn_o_1_381_0 = sub_353_d0;
  assign stage_0_sb = insn_o_1_381_0;
  assign insn_o_1_382_0 = stage_0_sb[15:0];
  assign stage_0_m0 = insn_o_1_382_0;
  assign insn_o_1_383_0 = stage_0_pr[15:0];
  assign stage_0_m1 = insn_o_1_383_0;
  assign insn_o_1_384_0 = stage_0_sb[16:16];
  assign stage_0_ms = insn_o_1_384_0;
  assign insn_o_1_385_0 = stage_0_ms ? stage_0_m1 : stage_0_m0;
  assign stage_0_mx = insn_o_1_385_0;
  assign insn_o_1_386_0 = zi_00[30:0];
  assign stage_0_zl = insn_o_1_386_0;
  assign insn_o_1_387_0 = ~stage_0_ms;
  assign stage_0_zb = insn_o_1_387_0;
  assign insn_o_1_388_0 = {stage_0_mx, stage_0_zl, stage_0_zb};
  assign stage_0_zo = insn_o_1_388_0;
  assign insn_o_1_389_0 = stage_0_zo[47:32];
  assign stage_0_zr = insn_o_1_389_0;
  assign insn_o_1_390_0 = stage_0_zo[31:0];
  assign stage_0_zq = insn_o_1_390_0;

  // Table 1
  always @(posedge clk) begin
    if (!rst_n) begin
      st_1_1 <= 0;
      st_1_2 <= 0;
      st_1_3 <= 0;
      st_1_4 <= 0;
      st_1_5 <= 0;
      st_1_6 <= 0;
      st_1_7 <= 0;
      st_1_8 <= 0;
      st_1_9 <= 0;
      st_1_10 <= 0;
      st_1_11 <= 0;
      st_1_12 <= 0;
      st_1_13 <= 0;
      st_1_14 <= 0;
      st_1_15 <= 0;
      st_1_16 <= 0;
      st_1_17 <= 0;
      st_1_18 <= 0;
      st_1_19 <= 0;
      st_1_20 <= 0;
      st_1_21 <= 0;
      st_1_22 <= 0;
      st_1_23 <= 0;
      st_1_24 <= 0;
      st_1_25 <= 0;
      st_1_26 <= 0;
      st_1_27 <= 0;
      st_1_28 <= 0;
      st_1_29 <= 0;
      st_1_30 <= 0;
      st_1_31 <= 0;
      st_1_32 <= 0;
      st_1_33 <= 0;
    end else begin
      if (start) begin
          zi_31 <= stage_32_zi_i;
          di_31 <= insn_o_1_6_0;
      end
      st_1_2 <= start;
      if (st_1_2) begin
          zi_30 <= stage_31_zo;
          di_30 <= di_31;
      end
      st_1_3 <= st_1_2;
      if (st_1_3) begin
          zi_29 <= stage_30_zo;
          di_29 <= di_30;
      end
      st_1_4 <= st_1_3;
      if (st_1_4) begin
          zi_28 <= stage_29_zo;
          di_28 <= di_29;
      end
      st_1_5 <= st_1_4;
      if (st_1_5) begin
          zi_27 <= stage_28_zo;
          di_27 <= di_28;
      end
      st_1_6 <= st_1_5;
      if (st_1_6) begin
          zi_26 <= stage_27_zo;
          di_26 <= di_27;
      end
      st_1_7 <= st_1_6;
      if (st_1_7) begin
          zi_25 <= stage_26_zo;
          di_25 <= di_26;
      end
      st_1_8 <= st_1_7;
      if (st_1_8) begin
          zi_24 <= stage_25_zo;
          di_24 <= di_25;
      end
      st_1_9 <= st_1_8;
      if (st_1_9) begin
          zi_23 <= stage_24_zo;
          di_23 <= di_24;
      end
      st_1_10 <= st_1_9;
      if (st_1_10) begin
          zi_22 <= stage_23_zo;
          di_22 <= di_23;
      end
      st_1_11 <= st_1_10;
      if (st_1_11) begin
          zi_21 <= stage_22_zo;
          di_21 <= di_22;
      end
      st_1_12 <= st_1_11;
      if (st_1_12) begin
          zi_20 <= stage_21_zo;
          di_20 <= di_21;
      end
      st_1_13 <= st_1_12;
      if (st_1_13) begin
          zi_19 <= stage_20_zo;
          di_19 <= di_20;
      end
      st_1_14 <= st_1_13;
      if (st_1_14) begin
          zi_18 <= stage_19_zo;
          di_18 <= di_19;
      end
      st_1_15 <= st_1_14;
      if (st_1_15) begin
          zi_17 <= stage_18_zo;
          di_17 <= di_18;
      end
      st_1_16 <= st_1_15;
      if (st_1_16) begin
          zi_16 <= stage_17_zo;
          di_16 <= di_17;
      end
      st_1_17 <= st_1_16;
      if (st_1_17) begin
          zi_15 <= stage_16_zo;
          di_15 <= di_16;
      end
      st_1_18 <= st_1_17;
      if (st_1_18) begin
          zi_14 <= stage_15_zo;
          di_14 <= di_15;
      end
      st_1_19 <= st_1_18;
      if (st_1_19) begin
          zi_13 <= stage_14_zo;
          di_13 <= di_14;
      end
      st_1_20 <= st_1_19;
      if (st_1_20) begin
          zi_12 <= stage_13_zo;
          di_12 <= di_13;
      end
      st_1_21 <= st_1_20;
      if (st_1_21) begin
          zi_11 <= stage_12_zo;
          di_11 <= di_12;
      end
      st_1_22 <= st_1_21;
      if (st_1_22) begin
          zi_10 <= stage_11_zo;
          di_10 <= di_11;
      end
      st_1_23 <= st_1_22;
      if (st_1_23) begin
          zi_09 <= stage_10_zo;
          di_09 <= di_10;
      end
      st_1_24 <= st_1_23;
      if (st_1_24) begin
          zi_08 <= stage_9_zo;
          di_08 <= di_09;
      end
      st_1_25 <= st_1_24;
      if (st_1_25) begin
          zi_07 <= stage_8_zo;
          di_07 <= di_08;
      end
      st_1_26 <= st_1_25;
      if (st_1_26) begin
          zi_06 <= stage_7_zo;
          di_06 <= di_07;
      end
      st_1_27 <= st_1_26;
      if (st_1_27) begin
          zi_05 <= stage_6_zo;
          di_05 <= di_06;
      end
      st_1_28 <= st_1_27;
      if (st_1_28) begin
          zi_04 <= stage_5_zo;
          di_04 <= di_05;
      end
      st_1_29 <= st_1_28;
      if (st_1_29) begin
          zi_03 <= stage_4_zo;
          di_03 <= di_04;
      end
      st_1_30 <= st_1_29;
      if (st_1_30) begin
          zi_02 <= stage_3_zo;
          di_02 <= di_03;
      end
      st_1_31 <= st_1_30;
      if (st_1_31) begin
          zi_01 <= stage_2_zo;
          di_01 <= di_02;
      end
      st_1_32 <= st_1_31;
      if (st_1_32) begin
          zi_00 <= stage_1_zo;
          di_00 <= di_01;
      end
      st_1_33 <= st_1_32;
      if (st_1_33) begin
          quotient <= stage_0_zq;
          remainder <= stage_0_zr;
      end
    end
  end

endmodule
