// Generated from iroha-0.1.0.

module fdiv(clk, rst_n, i_valid, z_out, z_valid, a_in, b_in);
  input clk;
  input rst_n;
  input i_valid;
  output [31:0] z_out;
  output z_valid;
  input [31:0] a_in;
  input [31:0] b_in;
  reg [31:0] z_out;
  reg z_valid;

  // State decls
  reg st_1_1;
  reg st_1_2;
  reg st_1_3;
  reg st_1_4;
  reg st_1_5;
  reg st_1_6;
  reg st_1_7;
  reg st_1_8;
  reg st_1_9;
  reg st_1_10;
  reg st_1_11;
  reg st_1_12;
  reg st_1_13;
  reg st_1_14;
  reg st_1_15;
  reg st_1_16;
  reg st_1_17;
  reg st_1_18;
  reg st_1_19;
  reg st_1_20;
  reg st_1_21;
  reg st_1_22;
  reg st_1_23;
  reg st_1_24;
  reg st_1_25;
  reg st_1_26;
  reg st_1_27;
  reg st_1_28;
  reg st_1_29;
  reg st_1_30;
  reg st_1_31;
  reg st_1_32;
  reg st_1_33;
  reg st_1_34;
  reg st_1_35;
  reg st_1_36;
  reg st_1_37;
  reg st_1_38;
  reg st_1_39;
  reg st_1_40;
  reg st_1_41;
  reg st_1_42;
  reg st_1_43;
  reg st_1_44;
  reg st_1_45;
  reg st_1_46;
  reg st_1_47;
  reg st_1_48;
  reg st_1_49;
  reg st_1_50;
  reg st_1_51;
  reg st_1_52;
  reg st_1_53;
  reg st_1_54;
  reg st_1_55;
  // State vars
  // Registers
  wire  [0:0] start;
  reg  [23:0] stage1_a_fraction;
  reg  [7:0] stage1_a_exponent;
  reg  stage1_a_sign;
  reg  stage1_a_exponent_is_all_0;
  reg  stage1_a_fraction_is_all_0;
  reg  [23:0] stage1_b_fraction;
  reg  [7:0] stage1_b_exponent;
  reg  stage1_b_sign;
  reg  stage1_b_exponent_is_all_0;
  reg  stage1_b_fraction_is_all_0;
  reg  [73:0] stage2_zi_00;
  reg  [73:0] stage2_zi_01;
  reg  [73:0] stage2_zi_02;
  reg  [73:0] stage2_zi_03;
  reg  [73:0] stage2_zi_04;
  reg  [73:0] stage2_zi_05;
  reg  [73:0] stage2_zi_06;
  reg  [73:0] stage2_zi_07;
  reg  [73:0] stage2_zi_08;
  reg  [73:0] stage2_zi_09;
  reg  [73:0] stage2_zi_10;
  reg  [73:0] stage2_zi_11;
  reg  [73:0] stage2_zi_12;
  reg  [73:0] stage2_zi_13;
  reg  [73:0] stage2_zi_14;
  reg  [73:0] stage2_zi_15;
  reg  [73:0] stage2_zi_16;
  reg  [73:0] stage2_zi_17;
  reg  [73:0] stage2_zi_18;
  reg  [73:0] stage2_zi_19;
  reg  [73:0] stage2_zi_20;
  reg  [73:0] stage2_zi_21;
  reg  [73:0] stage2_zi_22;
  reg  [73:0] stage2_zi_23;
  reg  [73:0] stage2_zi_24;
  reg  [73:0] stage2_zi_25;
  reg  [73:0] stage2_zi_26;
  reg  [73:0] stage2_zi_27;
  reg  [73:0] stage2_zi_28;
  reg  [73:0] stage2_zi_29;
  reg  [73:0] stage2_zi_30;
  reg  [73:0] stage2_zi_31;
  reg  [73:0] stage2_zi_32;
  reg  [73:0] stage2_zi_33;
  reg  [73:0] stage2_zi_34;
  reg  [73:0] stage2_zi_35;
  reg  [73:0] stage2_zi_36;
  reg  [73:0] stage2_zi_37;
  reg  [73:0] stage2_zi_38;
  reg  [73:0] stage2_zi_39;
  reg  [73:0] stage2_zi_40;
  reg  [73:0] stage2_zi_41;
  reg  [73:0] stage2_zi_42;
  reg  [73:0] stage2_zi_43;
  reg  [73:0] stage2_zi_44;
  reg  [73:0] stage2_zi_45;
  reg  [73:0] stage2_zi_46;
  reg  [73:0] stage2_zi_47;
  reg  [73:0] stage2_zi_48;
  reg  [73:0] stage2_zi_49;
  reg  [73:0] stage2_zi_50;
  reg  [23:0] stage2_di_00;
  reg  [23:0] stage2_di_01;
  reg  [23:0] stage2_di_02;
  reg  [23:0] stage2_di_03;
  reg  [23:0] stage2_di_04;
  reg  [23:0] stage2_di_05;
  reg  [23:0] stage2_di_06;
  reg  [23:0] stage2_di_07;
  reg  [23:0] stage2_di_08;
  reg  [23:0] stage2_di_09;
  reg  [23:0] stage2_di_10;
  reg  [23:0] stage2_di_11;
  reg  [23:0] stage2_di_12;
  reg  [23:0] stage2_di_13;
  reg  [23:0] stage2_di_14;
  reg  [23:0] stage2_di_15;
  reg  [23:0] stage2_di_16;
  reg  [23:0] stage2_di_17;
  reg  [23:0] stage2_di_18;
  reg  [23:0] stage2_di_19;
  reg  [23:0] stage2_di_20;
  reg  [23:0] stage2_di_21;
  reg  [23:0] stage2_di_22;
  reg  [23:0] stage2_di_23;
  reg  [23:0] stage2_di_24;
  reg  [23:0] stage2_di_25;
  reg  [23:0] stage2_di_26;
  reg  [23:0] stage2_di_27;
  reg  [23:0] stage2_di_28;
  reg  [23:0] stage2_di_29;
  reg  [23:0] stage2_di_30;
  reg  [23:0] stage2_di_31;
  reg  [23:0] stage2_di_32;
  reg  [23:0] stage2_di_33;
  reg  [23:0] stage2_di_34;
  reg  [23:0] stage2_di_35;
  reg  [23:0] stage2_di_36;
  reg  [23:0] stage2_di_37;
  reg  [23:0] stage2_di_38;
  reg  [23:0] stage2_di_39;
  reg  [23:0] stage2_di_40;
  reg  [23:0] stage2_di_41;
  reg  [23:0] stage2_di_42;
  reg  [23:0] stage2_di_43;
  reg  [23:0] stage2_di_44;
  reg  [23:0] stage2_di_45;
  reg  [23:0] stage2_di_46;
  reg  [23:0] stage2_di_47;
  reg  [23:0] stage2_di_48;
  reg  [23:0] stage2_di_49;
  reg  [23:0] stage2_di_50;
  reg  signed [9:0] stage2_exponent_00;
  reg  signed [9:0] stage2_exponent_01;
  reg  signed [9:0] stage2_exponent_02;
  reg  signed [9:0] stage2_exponent_03;
  reg  signed [9:0] stage2_exponent_04;
  reg  signed [9:0] stage2_exponent_05;
  reg  signed [9:0] stage2_exponent_06;
  reg  signed [9:0] stage2_exponent_07;
  reg  signed [9:0] stage2_exponent_08;
  reg  signed [9:0] stage2_exponent_09;
  reg  signed [9:0] stage2_exponent_10;
  reg  signed [9:0] stage2_exponent_11;
  reg  signed [9:0] stage2_exponent_12;
  reg  signed [9:0] stage2_exponent_13;
  reg  signed [9:0] stage2_exponent_14;
  reg  signed [9:0] stage2_exponent_15;
  reg  signed [9:0] stage2_exponent_16;
  reg  signed [9:0] stage2_exponent_17;
  reg  signed [9:0] stage2_exponent_18;
  reg  signed [9:0] stage2_exponent_19;
  reg  signed [9:0] stage2_exponent_20;
  reg  signed [9:0] stage2_exponent_21;
  reg  signed [9:0] stage2_exponent_22;
  reg  signed [9:0] stage2_exponent_23;
  reg  signed [9:0] stage2_exponent_24;
  reg  signed [9:0] stage2_exponent_25;
  reg  signed [9:0] stage2_exponent_26;
  reg  signed [9:0] stage2_exponent_27;
  reg  signed [9:0] stage2_exponent_28;
  reg  signed [9:0] stage2_exponent_29;
  reg  signed [9:0] stage2_exponent_30;
  reg  signed [9:0] stage2_exponent_31;
  reg  signed [9:0] stage2_exponent_32;
  reg  signed [9:0] stage2_exponent_33;
  reg  signed [9:0] stage2_exponent_34;
  reg  signed [9:0] stage2_exponent_35;
  reg  signed [9:0] stage2_exponent_36;
  reg  signed [9:0] stage2_exponent_37;
  reg  signed [9:0] stage2_exponent_38;
  reg  signed [9:0] stage2_exponent_39;
  reg  signed [9:0] stage2_exponent_40;
  reg  signed [9:0] stage2_exponent_41;
  reg  signed [9:0] stage2_exponent_42;
  reg  signed [9:0] stage2_exponent_43;
  reg  signed [9:0] stage2_exponent_44;
  reg  signed [9:0] stage2_exponent_45;
  reg  signed [9:0] stage2_exponent_46;
  reg  signed [9:0] stage2_exponent_47;
  reg  signed [9:0] stage2_exponent_48;
  reg  signed [9:0] stage2_exponent_49;
  reg  signed [9:0] stage2_exponent_50;
  reg  stage2_sign_00;
  reg  stage2_sign_01;
  reg  stage2_sign_02;
  reg  stage2_sign_03;
  reg  stage2_sign_04;
  reg  stage2_sign_05;
  reg  stage2_sign_06;
  reg  stage2_sign_07;
  reg  stage2_sign_08;
  reg  stage2_sign_09;
  reg  stage2_sign_10;
  reg  stage2_sign_11;
  reg  stage2_sign_12;
  reg  stage2_sign_13;
  reg  stage2_sign_14;
  reg  stage2_sign_15;
  reg  stage2_sign_16;
  reg  stage2_sign_17;
  reg  stage2_sign_18;
  reg  stage2_sign_19;
  reg  stage2_sign_20;
  reg  stage2_sign_21;
  reg  stage2_sign_22;
  reg  stage2_sign_23;
  reg  stage2_sign_24;
  reg  stage2_sign_25;
  reg  stage2_sign_26;
  reg  stage2_sign_27;
  reg  stage2_sign_28;
  reg  stage2_sign_29;
  reg  stage2_sign_30;
  reg  stage2_sign_31;
  reg  stage2_sign_32;
  reg  stage2_sign_33;
  reg  stage2_sign_34;
  reg  stage2_sign_35;
  reg  stage2_sign_36;
  reg  stage2_sign_37;
  reg  stage2_sign_38;
  reg  stage2_sign_39;
  reg  stage2_sign_40;
  reg  stage2_sign_41;
  reg  stage2_sign_42;
  reg  stage2_sign_43;
  reg  stage2_sign_44;
  reg  stage2_sign_45;
  reg  stage2_sign_46;
  reg  stage2_sign_47;
  reg  stage2_sign_48;
  reg  stage2_sign_49;
  reg  stage2_sign_50;
  reg  stage2_a_is_zero_00;
  reg  stage2_a_is_zero_01;
  reg  stage2_a_is_zero_02;
  reg  stage2_a_is_zero_03;
  reg  stage2_a_is_zero_04;
  reg  stage2_a_is_zero_05;
  reg  stage2_a_is_zero_06;
  reg  stage2_a_is_zero_07;
  reg  stage2_a_is_zero_08;
  reg  stage2_a_is_zero_09;
  reg  stage2_a_is_zero_10;
  reg  stage2_a_is_zero_11;
  reg  stage2_a_is_zero_12;
  reg  stage2_a_is_zero_13;
  reg  stage2_a_is_zero_14;
  reg  stage2_a_is_zero_15;
  reg  stage2_a_is_zero_16;
  reg  stage2_a_is_zero_17;
  reg  stage2_a_is_zero_18;
  reg  stage2_a_is_zero_19;
  reg  stage2_a_is_zero_20;
  reg  stage2_a_is_zero_21;
  reg  stage2_a_is_zero_22;
  reg  stage2_a_is_zero_23;
  reg  stage2_a_is_zero_24;
  reg  stage2_a_is_zero_25;
  reg  stage2_a_is_zero_26;
  reg  stage2_a_is_zero_27;
  reg  stage2_a_is_zero_28;
  reg  stage2_a_is_zero_29;
  reg  stage2_a_is_zero_30;
  reg  stage2_a_is_zero_31;
  reg  stage2_a_is_zero_32;
  reg  stage2_a_is_zero_33;
  reg  stage2_a_is_zero_34;
  reg  stage2_a_is_zero_35;
  reg  stage2_a_is_zero_36;
  reg  stage2_a_is_zero_37;
  reg  stage2_a_is_zero_38;
  reg  stage2_a_is_zero_39;
  reg  stage2_a_is_zero_40;
  reg  stage2_a_is_zero_41;
  reg  stage2_a_is_zero_42;
  reg  stage2_a_is_zero_43;
  reg  stage2_a_is_zero_44;
  reg  stage2_a_is_zero_45;
  reg  stage2_a_is_zero_46;
  reg  stage2_a_is_zero_47;
  reg  stage2_a_is_zero_48;
  reg  stage2_a_is_zero_49;
  reg  stage2_a_is_zero_50;
  reg  stage2_a_is_inf_00;
  reg  stage2_a_is_inf_01;
  reg  stage2_a_is_inf_02;
  reg  stage2_a_is_inf_03;
  reg  stage2_a_is_inf_04;
  reg  stage2_a_is_inf_05;
  reg  stage2_a_is_inf_06;
  reg  stage2_a_is_inf_07;
  reg  stage2_a_is_inf_08;
  reg  stage2_a_is_inf_09;
  reg  stage2_a_is_inf_10;
  reg  stage2_a_is_inf_11;
  reg  stage2_a_is_inf_12;
  reg  stage2_a_is_inf_13;
  reg  stage2_a_is_inf_14;
  reg  stage2_a_is_inf_15;
  reg  stage2_a_is_inf_16;
  reg  stage2_a_is_inf_17;
  reg  stage2_a_is_inf_18;
  reg  stage2_a_is_inf_19;
  reg  stage2_a_is_inf_20;
  reg  stage2_a_is_inf_21;
  reg  stage2_a_is_inf_22;
  reg  stage2_a_is_inf_23;
  reg  stage2_a_is_inf_24;
  reg  stage2_a_is_inf_25;
  reg  stage2_a_is_inf_26;
  reg  stage2_a_is_inf_27;
  reg  stage2_a_is_inf_28;
  reg  stage2_a_is_inf_29;
  reg  stage2_a_is_inf_30;
  reg  stage2_a_is_inf_31;
  reg  stage2_a_is_inf_32;
  reg  stage2_a_is_inf_33;
  reg  stage2_a_is_inf_34;
  reg  stage2_a_is_inf_35;
  reg  stage2_a_is_inf_36;
  reg  stage2_a_is_inf_37;
  reg  stage2_a_is_inf_38;
  reg  stage2_a_is_inf_39;
  reg  stage2_a_is_inf_40;
  reg  stage2_a_is_inf_41;
  reg  stage2_a_is_inf_42;
  reg  stage2_a_is_inf_43;
  reg  stage2_a_is_inf_44;
  reg  stage2_a_is_inf_45;
  reg  stage2_a_is_inf_46;
  reg  stage2_a_is_inf_47;
  reg  stage2_a_is_inf_48;
  reg  stage2_a_is_inf_49;
  reg  stage2_a_is_inf_50;
  reg  stage2_a_is_nan_00;
  reg  stage2_a_is_nan_01;
  reg  stage2_a_is_nan_02;
  reg  stage2_a_is_nan_03;
  reg  stage2_a_is_nan_04;
  reg  stage2_a_is_nan_05;
  reg  stage2_a_is_nan_06;
  reg  stage2_a_is_nan_07;
  reg  stage2_a_is_nan_08;
  reg  stage2_a_is_nan_09;
  reg  stage2_a_is_nan_10;
  reg  stage2_a_is_nan_11;
  reg  stage2_a_is_nan_12;
  reg  stage2_a_is_nan_13;
  reg  stage2_a_is_nan_14;
  reg  stage2_a_is_nan_15;
  reg  stage2_a_is_nan_16;
  reg  stage2_a_is_nan_17;
  reg  stage2_a_is_nan_18;
  reg  stage2_a_is_nan_19;
  reg  stage2_a_is_nan_20;
  reg  stage2_a_is_nan_21;
  reg  stage2_a_is_nan_22;
  reg  stage2_a_is_nan_23;
  reg  stage2_a_is_nan_24;
  reg  stage2_a_is_nan_25;
  reg  stage2_a_is_nan_26;
  reg  stage2_a_is_nan_27;
  reg  stage2_a_is_nan_28;
  reg  stage2_a_is_nan_29;
  reg  stage2_a_is_nan_30;
  reg  stage2_a_is_nan_31;
  reg  stage2_a_is_nan_32;
  reg  stage2_a_is_nan_33;
  reg  stage2_a_is_nan_34;
  reg  stage2_a_is_nan_35;
  reg  stage2_a_is_nan_36;
  reg  stage2_a_is_nan_37;
  reg  stage2_a_is_nan_38;
  reg  stage2_a_is_nan_39;
  reg  stage2_a_is_nan_40;
  reg  stage2_a_is_nan_41;
  reg  stage2_a_is_nan_42;
  reg  stage2_a_is_nan_43;
  reg  stage2_a_is_nan_44;
  reg  stage2_a_is_nan_45;
  reg  stage2_a_is_nan_46;
  reg  stage2_a_is_nan_47;
  reg  stage2_a_is_nan_48;
  reg  stage2_a_is_nan_49;
  reg  stage2_a_is_nan_50;
  reg  stage2_b_is_zero_00;
  reg  stage2_b_is_zero_01;
  reg  stage2_b_is_zero_02;
  reg  stage2_b_is_zero_03;
  reg  stage2_b_is_zero_04;
  reg  stage2_b_is_zero_05;
  reg  stage2_b_is_zero_06;
  reg  stage2_b_is_zero_07;
  reg  stage2_b_is_zero_08;
  reg  stage2_b_is_zero_09;
  reg  stage2_b_is_zero_10;
  reg  stage2_b_is_zero_11;
  reg  stage2_b_is_zero_12;
  reg  stage2_b_is_zero_13;
  reg  stage2_b_is_zero_14;
  reg  stage2_b_is_zero_15;
  reg  stage2_b_is_zero_16;
  reg  stage2_b_is_zero_17;
  reg  stage2_b_is_zero_18;
  reg  stage2_b_is_zero_19;
  reg  stage2_b_is_zero_20;
  reg  stage2_b_is_zero_21;
  reg  stage2_b_is_zero_22;
  reg  stage2_b_is_zero_23;
  reg  stage2_b_is_zero_24;
  reg  stage2_b_is_zero_25;
  reg  stage2_b_is_zero_26;
  reg  stage2_b_is_zero_27;
  reg  stage2_b_is_zero_28;
  reg  stage2_b_is_zero_29;
  reg  stage2_b_is_zero_30;
  reg  stage2_b_is_zero_31;
  reg  stage2_b_is_zero_32;
  reg  stage2_b_is_zero_33;
  reg  stage2_b_is_zero_34;
  reg  stage2_b_is_zero_35;
  reg  stage2_b_is_zero_36;
  reg  stage2_b_is_zero_37;
  reg  stage2_b_is_zero_38;
  reg  stage2_b_is_zero_39;
  reg  stage2_b_is_zero_40;
  reg  stage2_b_is_zero_41;
  reg  stage2_b_is_zero_42;
  reg  stage2_b_is_zero_43;
  reg  stage2_b_is_zero_44;
  reg  stage2_b_is_zero_45;
  reg  stage2_b_is_zero_46;
  reg  stage2_b_is_zero_47;
  reg  stage2_b_is_zero_48;
  reg  stage2_b_is_zero_49;
  reg  stage2_b_is_zero_50;
  reg  stage2_b_is_inf_00;
  reg  stage2_b_is_inf_01;
  reg  stage2_b_is_inf_02;
  reg  stage2_b_is_inf_03;
  reg  stage2_b_is_inf_04;
  reg  stage2_b_is_inf_05;
  reg  stage2_b_is_inf_06;
  reg  stage2_b_is_inf_07;
  reg  stage2_b_is_inf_08;
  reg  stage2_b_is_inf_09;
  reg  stage2_b_is_inf_10;
  reg  stage2_b_is_inf_11;
  reg  stage2_b_is_inf_12;
  reg  stage2_b_is_inf_13;
  reg  stage2_b_is_inf_14;
  reg  stage2_b_is_inf_15;
  reg  stage2_b_is_inf_16;
  reg  stage2_b_is_inf_17;
  reg  stage2_b_is_inf_18;
  reg  stage2_b_is_inf_19;
  reg  stage2_b_is_inf_20;
  reg  stage2_b_is_inf_21;
  reg  stage2_b_is_inf_22;
  reg  stage2_b_is_inf_23;
  reg  stage2_b_is_inf_24;
  reg  stage2_b_is_inf_25;
  reg  stage2_b_is_inf_26;
  reg  stage2_b_is_inf_27;
  reg  stage2_b_is_inf_28;
  reg  stage2_b_is_inf_29;
  reg  stage2_b_is_inf_30;
  reg  stage2_b_is_inf_31;
  reg  stage2_b_is_inf_32;
  reg  stage2_b_is_inf_33;
  reg  stage2_b_is_inf_34;
  reg  stage2_b_is_inf_35;
  reg  stage2_b_is_inf_36;
  reg  stage2_b_is_inf_37;
  reg  stage2_b_is_inf_38;
  reg  stage2_b_is_inf_39;
  reg  stage2_b_is_inf_40;
  reg  stage2_b_is_inf_41;
  reg  stage2_b_is_inf_42;
  reg  stage2_b_is_inf_43;
  reg  stage2_b_is_inf_44;
  reg  stage2_b_is_inf_45;
  reg  stage2_b_is_inf_46;
  reg  stage2_b_is_inf_47;
  reg  stage2_b_is_inf_48;
  reg  stage2_b_is_inf_49;
  reg  stage2_b_is_inf_50;
  reg  stage2_b_is_nan_00;
  reg  stage2_b_is_nan_01;
  reg  stage2_b_is_nan_02;
  reg  stage2_b_is_nan_03;
  reg  stage2_b_is_nan_04;
  reg  stage2_b_is_nan_05;
  reg  stage2_b_is_nan_06;
  reg  stage2_b_is_nan_07;
  reg  stage2_b_is_nan_08;
  reg  stage2_b_is_nan_09;
  reg  stage2_b_is_nan_10;
  reg  stage2_b_is_nan_11;
  reg  stage2_b_is_nan_12;
  reg  stage2_b_is_nan_13;
  reg  stage2_b_is_nan_14;
  reg  stage2_b_is_nan_15;
  reg  stage2_b_is_nan_16;
  reg  stage2_b_is_nan_17;
  reg  stage2_b_is_nan_18;
  reg  stage2_b_is_nan_19;
  reg  stage2_b_is_nan_20;
  reg  stage2_b_is_nan_21;
  reg  stage2_b_is_nan_22;
  reg  stage2_b_is_nan_23;
  reg  stage2_b_is_nan_24;
  reg  stage2_b_is_nan_25;
  reg  stage2_b_is_nan_26;
  reg  stage2_b_is_nan_27;
  reg  stage2_b_is_nan_28;
  reg  stage2_b_is_nan_29;
  reg  stage2_b_is_nan_30;
  reg  stage2_b_is_nan_31;
  reg  stage2_b_is_nan_32;
  reg  stage2_b_is_nan_33;
  reg  stage2_b_is_nan_34;
  reg  stage2_b_is_nan_35;
  reg  stage2_b_is_nan_36;
  reg  stage2_b_is_nan_37;
  reg  stage2_b_is_nan_38;
  reg  stage2_b_is_nan_39;
  reg  stage2_b_is_nan_40;
  reg  stage2_b_is_nan_41;
  reg  stage2_b_is_nan_42;
  reg  stage2_b_is_nan_43;
  reg  stage2_b_is_nan_44;
  reg  stage2_b_is_nan_45;
  reg  stage2_b_is_nan_46;
  reg  stage2_b_is_nan_47;
  reg  stage2_b_is_nan_48;
  reg  stage2_b_is_nan_49;
  reg  stage2_b_is_nan_50;
  reg  [26:0] stage3_fraction;
  reg  signed [9:0] stage3_exponent;
  reg  stage3_sign;
  reg  stage3_a_is_zero;
  reg  stage3_a_is_inf;
  reg  stage3_a_is_nan;
  reg  stage3_b_is_zero;
  reg  stage3_b_is_inf;
  reg  stage3_b_is_nan;
  reg  [23:0] stage4_fraction;
  reg  signed [9:0] stage4_exponent;
  reg  stage4_sign;
  reg  stage4_a_is_zero;
  reg  stage4_a_is_inf;
  reg  stage4_a_is_nan;
  reg  stage4_b_is_zero;
  reg  stage4_b_is_inf;
  reg  stage4_b_is_nan;
  wire  [31:0] stage1_a_data_in;
  wire  [7:0] stage1_a_exponent_in;
  wire  [22:0] stage1_a_fraction_in;
  wire  stage1_a_sign_in;
  wire  stage1_a_exponent_zero;
  wire  [0:0] stage1_a_fraction_msb;
  wire  [31:0] stage1_b_data_in;
  wire  [7:0] stage1_b_exponent_in;
  wire  [22:0] stage1_b_fraction_in;
  wire  stage1_b_sign_in;
  wire  stage1_b_exponent_zero;
  wire  [0:0] stage1_b_fraction_msb;
  wire  [9:0] stage2_50_exponent_a_in;
  wire  signed [9:0] stage2_50_exponent_a_d;
  wire  [9:0] stage2_50_exponent_b_in;
  wire  signed [9:0] stage2_50_exponent_b_d;
  wire  stage2_50_exponent_a_is_all_0;
  wire  stage2_50_exponent_a_is_all_1;
  wire  stage2_50_fraction_a_is_all_0;
  wire  stage2_50_fraction_a_is_not_0;
  wire  stage2_50_exponent_b_is_all_0;
  wire  stage2_50_exponent_b_is_all_1;
  wire  stage2_50_fraction_b_is_all_0;
  wire  stage2_50_fraction_b_is_not_0;
  wire  [24:0] stage2_49_pr;
  wire  [24:0] stage2_49_sb;
  wire  [23:0] stage2_49_m0;
  wire  [23:0] stage2_49_m1;
  wire  [0:0] stage2_49_ms;
  wire  [23:0] stage2_49_mx;
  wire  [48:0] stage2_49_zl;
  wire  [0:0] stage2_49_zb;
  wire  [24:0] stage2_48_pr;
  wire  [24:0] stage2_48_sb;
  wire  [23:0] stage2_48_m0;
  wire  [23:0] stage2_48_m1;
  wire  [0:0] stage2_48_ms;
  wire  [23:0] stage2_48_mx;
  wire  [48:0] stage2_48_zl;
  wire  [0:0] stage2_48_zb;
  wire  [24:0] stage2_47_pr;
  wire  [24:0] stage2_47_sb;
  wire  [23:0] stage2_47_m0;
  wire  [23:0] stage2_47_m1;
  wire  [0:0] stage2_47_ms;
  wire  [23:0] stage2_47_mx;
  wire  [48:0] stage2_47_zl;
  wire  [0:0] stage2_47_zb;
  wire  [24:0] stage2_46_pr;
  wire  [24:0] stage2_46_sb;
  wire  [23:0] stage2_46_m0;
  wire  [23:0] stage2_46_m1;
  wire  [0:0] stage2_46_ms;
  wire  [23:0] stage2_46_mx;
  wire  [48:0] stage2_46_zl;
  wire  [0:0] stage2_46_zb;
  wire  [24:0] stage2_45_pr;
  wire  [24:0] stage2_45_sb;
  wire  [23:0] stage2_45_m0;
  wire  [23:0] stage2_45_m1;
  wire  [0:0] stage2_45_ms;
  wire  [23:0] stage2_45_mx;
  wire  [48:0] stage2_45_zl;
  wire  [0:0] stage2_45_zb;
  wire  [24:0] stage2_44_pr;
  wire  [24:0] stage2_44_sb;
  wire  [23:0] stage2_44_m0;
  wire  [23:0] stage2_44_m1;
  wire  [0:0] stage2_44_ms;
  wire  [23:0] stage2_44_mx;
  wire  [48:0] stage2_44_zl;
  wire  [0:0] stage2_44_zb;
  wire  [24:0] stage2_43_pr;
  wire  [24:0] stage2_43_sb;
  wire  [23:0] stage2_43_m0;
  wire  [23:0] stage2_43_m1;
  wire  [0:0] stage2_43_ms;
  wire  [23:0] stage2_43_mx;
  wire  [48:0] stage2_43_zl;
  wire  [0:0] stage2_43_zb;
  wire  [24:0] stage2_42_pr;
  wire  [24:0] stage2_42_sb;
  wire  [23:0] stage2_42_m0;
  wire  [23:0] stage2_42_m1;
  wire  [0:0] stage2_42_ms;
  wire  [23:0] stage2_42_mx;
  wire  [48:0] stage2_42_zl;
  wire  [0:0] stage2_42_zb;
  wire  [24:0] stage2_41_pr;
  wire  [24:0] stage2_41_sb;
  wire  [23:0] stage2_41_m0;
  wire  [23:0] stage2_41_m1;
  wire  [0:0] stage2_41_ms;
  wire  [23:0] stage2_41_mx;
  wire  [48:0] stage2_41_zl;
  wire  [0:0] stage2_41_zb;
  wire  [24:0] stage2_40_pr;
  wire  [24:0] stage2_40_sb;
  wire  [23:0] stage2_40_m0;
  wire  [23:0] stage2_40_m1;
  wire  [0:0] stage2_40_ms;
  wire  [23:0] stage2_40_mx;
  wire  [48:0] stage2_40_zl;
  wire  [0:0] stage2_40_zb;
  wire  [24:0] stage2_39_pr;
  wire  [24:0] stage2_39_sb;
  wire  [23:0] stage2_39_m0;
  wire  [23:0] stage2_39_m1;
  wire  [0:0] stage2_39_ms;
  wire  [23:0] stage2_39_mx;
  wire  [48:0] stage2_39_zl;
  wire  [0:0] stage2_39_zb;
  wire  [24:0] stage2_38_pr;
  wire  [24:0] stage2_38_sb;
  wire  [23:0] stage2_38_m0;
  wire  [23:0] stage2_38_m1;
  wire  [0:0] stage2_38_ms;
  wire  [23:0] stage2_38_mx;
  wire  [48:0] stage2_38_zl;
  wire  [0:0] stage2_38_zb;
  wire  [24:0] stage2_37_pr;
  wire  [24:0] stage2_37_sb;
  wire  [23:0] stage2_37_m0;
  wire  [23:0] stage2_37_m1;
  wire  [0:0] stage2_37_ms;
  wire  [23:0] stage2_37_mx;
  wire  [48:0] stage2_37_zl;
  wire  [0:0] stage2_37_zb;
  wire  [24:0] stage2_36_pr;
  wire  [24:0] stage2_36_sb;
  wire  [23:0] stage2_36_m0;
  wire  [23:0] stage2_36_m1;
  wire  [0:0] stage2_36_ms;
  wire  [23:0] stage2_36_mx;
  wire  [48:0] stage2_36_zl;
  wire  [0:0] stage2_36_zb;
  wire  [24:0] stage2_35_pr;
  wire  [24:0] stage2_35_sb;
  wire  [23:0] stage2_35_m0;
  wire  [23:0] stage2_35_m1;
  wire  [0:0] stage2_35_ms;
  wire  [23:0] stage2_35_mx;
  wire  [48:0] stage2_35_zl;
  wire  [0:0] stage2_35_zb;
  wire  [24:0] stage2_34_pr;
  wire  [24:0] stage2_34_sb;
  wire  [23:0] stage2_34_m0;
  wire  [23:0] stage2_34_m1;
  wire  [0:0] stage2_34_ms;
  wire  [23:0] stage2_34_mx;
  wire  [48:0] stage2_34_zl;
  wire  [0:0] stage2_34_zb;
  wire  [24:0] stage2_33_pr;
  wire  [24:0] stage2_33_sb;
  wire  [23:0] stage2_33_m0;
  wire  [23:0] stage2_33_m1;
  wire  [0:0] stage2_33_ms;
  wire  [23:0] stage2_33_mx;
  wire  [48:0] stage2_33_zl;
  wire  [0:0] stage2_33_zb;
  wire  [24:0] stage2_32_pr;
  wire  [24:0] stage2_32_sb;
  wire  [23:0] stage2_32_m0;
  wire  [23:0] stage2_32_m1;
  wire  [0:0] stage2_32_ms;
  wire  [23:0] stage2_32_mx;
  wire  [48:0] stage2_32_zl;
  wire  [0:0] stage2_32_zb;
  wire  [24:0] stage2_31_pr;
  wire  [24:0] stage2_31_sb;
  wire  [23:0] stage2_31_m0;
  wire  [23:0] stage2_31_m1;
  wire  [0:0] stage2_31_ms;
  wire  [23:0] stage2_31_mx;
  wire  [48:0] stage2_31_zl;
  wire  [0:0] stage2_31_zb;
  wire  [24:0] stage2_30_pr;
  wire  [24:0] stage2_30_sb;
  wire  [23:0] stage2_30_m0;
  wire  [23:0] stage2_30_m1;
  wire  [0:0] stage2_30_ms;
  wire  [23:0] stage2_30_mx;
  wire  [48:0] stage2_30_zl;
  wire  [0:0] stage2_30_zb;
  wire  [24:0] stage2_29_pr;
  wire  [24:0] stage2_29_sb;
  wire  [23:0] stage2_29_m0;
  wire  [23:0] stage2_29_m1;
  wire  [0:0] stage2_29_ms;
  wire  [23:0] stage2_29_mx;
  wire  [48:0] stage2_29_zl;
  wire  [0:0] stage2_29_zb;
  wire  [24:0] stage2_28_pr;
  wire  [24:0] stage2_28_sb;
  wire  [23:0] stage2_28_m0;
  wire  [23:0] stage2_28_m1;
  wire  [0:0] stage2_28_ms;
  wire  [23:0] stage2_28_mx;
  wire  [48:0] stage2_28_zl;
  wire  [0:0] stage2_28_zb;
  wire  [24:0] stage2_27_pr;
  wire  [24:0] stage2_27_sb;
  wire  [23:0] stage2_27_m0;
  wire  [23:0] stage2_27_m1;
  wire  [0:0] stage2_27_ms;
  wire  [23:0] stage2_27_mx;
  wire  [48:0] stage2_27_zl;
  wire  [0:0] stage2_27_zb;
  wire  [24:0] stage2_26_pr;
  wire  [24:0] stage2_26_sb;
  wire  [23:0] stage2_26_m0;
  wire  [23:0] stage2_26_m1;
  wire  [0:0] stage2_26_ms;
  wire  [23:0] stage2_26_mx;
  wire  [48:0] stage2_26_zl;
  wire  [0:0] stage2_26_zb;
  wire  [24:0] stage2_25_pr;
  wire  [24:0] stage2_25_sb;
  wire  [23:0] stage2_25_m0;
  wire  [23:0] stage2_25_m1;
  wire  [0:0] stage2_25_ms;
  wire  [23:0] stage2_25_mx;
  wire  [48:0] stage2_25_zl;
  wire  [0:0] stage2_25_zb;
  wire  [24:0] stage2_24_pr;
  wire  [24:0] stage2_24_sb;
  wire  [23:0] stage2_24_m0;
  wire  [23:0] stage2_24_m1;
  wire  [0:0] stage2_24_ms;
  wire  [23:0] stage2_24_mx;
  wire  [48:0] stage2_24_zl;
  wire  [0:0] stage2_24_zb;
  wire  [24:0] stage2_23_pr;
  wire  [24:0] stage2_23_sb;
  wire  [23:0] stage2_23_m0;
  wire  [23:0] stage2_23_m1;
  wire  [0:0] stage2_23_ms;
  wire  [23:0] stage2_23_mx;
  wire  [48:0] stage2_23_zl;
  wire  [0:0] stage2_23_zb;
  wire  [24:0] stage2_22_pr;
  wire  [24:0] stage2_22_sb;
  wire  [23:0] stage2_22_m0;
  wire  [23:0] stage2_22_m1;
  wire  [0:0] stage2_22_ms;
  wire  [23:0] stage2_22_mx;
  wire  [48:0] stage2_22_zl;
  wire  [0:0] stage2_22_zb;
  wire  [24:0] stage2_21_pr;
  wire  [24:0] stage2_21_sb;
  wire  [23:0] stage2_21_m0;
  wire  [23:0] stage2_21_m1;
  wire  [0:0] stage2_21_ms;
  wire  [23:0] stage2_21_mx;
  wire  [48:0] stage2_21_zl;
  wire  [0:0] stage2_21_zb;
  wire  [24:0] stage2_20_pr;
  wire  [24:0] stage2_20_sb;
  wire  [23:0] stage2_20_m0;
  wire  [23:0] stage2_20_m1;
  wire  [0:0] stage2_20_ms;
  wire  [23:0] stage2_20_mx;
  wire  [48:0] stage2_20_zl;
  wire  [0:0] stage2_20_zb;
  wire  [24:0] stage2_19_pr;
  wire  [24:0] stage2_19_sb;
  wire  [23:0] stage2_19_m0;
  wire  [23:0] stage2_19_m1;
  wire  [0:0] stage2_19_ms;
  wire  [23:0] stage2_19_mx;
  wire  [48:0] stage2_19_zl;
  wire  [0:0] stage2_19_zb;
  wire  [24:0] stage2_18_pr;
  wire  [24:0] stage2_18_sb;
  wire  [23:0] stage2_18_m0;
  wire  [23:0] stage2_18_m1;
  wire  [0:0] stage2_18_ms;
  wire  [23:0] stage2_18_mx;
  wire  [48:0] stage2_18_zl;
  wire  [0:0] stage2_18_zb;
  wire  [24:0] stage2_17_pr;
  wire  [24:0] stage2_17_sb;
  wire  [23:0] stage2_17_m0;
  wire  [23:0] stage2_17_m1;
  wire  [0:0] stage2_17_ms;
  wire  [23:0] stage2_17_mx;
  wire  [48:0] stage2_17_zl;
  wire  [0:0] stage2_17_zb;
  wire  [24:0] stage2_16_pr;
  wire  [24:0] stage2_16_sb;
  wire  [23:0] stage2_16_m0;
  wire  [23:0] stage2_16_m1;
  wire  [0:0] stage2_16_ms;
  wire  [23:0] stage2_16_mx;
  wire  [48:0] stage2_16_zl;
  wire  [0:0] stage2_16_zb;
  wire  [24:0] stage2_15_pr;
  wire  [24:0] stage2_15_sb;
  wire  [23:0] stage2_15_m0;
  wire  [23:0] stage2_15_m1;
  wire  [0:0] stage2_15_ms;
  wire  [23:0] stage2_15_mx;
  wire  [48:0] stage2_15_zl;
  wire  [0:0] stage2_15_zb;
  wire  [24:0] stage2_14_pr;
  wire  [24:0] stage2_14_sb;
  wire  [23:0] stage2_14_m0;
  wire  [23:0] stage2_14_m1;
  wire  [0:0] stage2_14_ms;
  wire  [23:0] stage2_14_mx;
  wire  [48:0] stage2_14_zl;
  wire  [0:0] stage2_14_zb;
  wire  [24:0] stage2_13_pr;
  wire  [24:0] stage2_13_sb;
  wire  [23:0] stage2_13_m0;
  wire  [23:0] stage2_13_m1;
  wire  [0:0] stage2_13_ms;
  wire  [23:0] stage2_13_mx;
  wire  [48:0] stage2_13_zl;
  wire  [0:0] stage2_13_zb;
  wire  [24:0] stage2_12_pr;
  wire  [24:0] stage2_12_sb;
  wire  [23:0] stage2_12_m0;
  wire  [23:0] stage2_12_m1;
  wire  [0:0] stage2_12_ms;
  wire  [23:0] stage2_12_mx;
  wire  [48:0] stage2_12_zl;
  wire  [0:0] stage2_12_zb;
  wire  [24:0] stage2_11_pr;
  wire  [24:0] stage2_11_sb;
  wire  [23:0] stage2_11_m0;
  wire  [23:0] stage2_11_m1;
  wire  [0:0] stage2_11_ms;
  wire  [23:0] stage2_11_mx;
  wire  [48:0] stage2_11_zl;
  wire  [0:0] stage2_11_zb;
  wire  [24:0] stage2_10_pr;
  wire  [24:0] stage2_10_sb;
  wire  [23:0] stage2_10_m0;
  wire  [23:0] stage2_10_m1;
  wire  [0:0] stage2_10_ms;
  wire  [23:0] stage2_10_mx;
  wire  [48:0] stage2_10_zl;
  wire  [0:0] stage2_10_zb;
  wire  [24:0] stage2_9_pr;
  wire  [24:0] stage2_9_sb;
  wire  [23:0] stage2_9_m0;
  wire  [23:0] stage2_9_m1;
  wire  [0:0] stage2_9_ms;
  wire  [23:0] stage2_9_mx;
  wire  [48:0] stage2_9_zl;
  wire  [0:0] stage2_9_zb;
  wire  [24:0] stage2_8_pr;
  wire  [24:0] stage2_8_sb;
  wire  [23:0] stage2_8_m0;
  wire  [23:0] stage2_8_m1;
  wire  [0:0] stage2_8_ms;
  wire  [23:0] stage2_8_mx;
  wire  [48:0] stage2_8_zl;
  wire  [0:0] stage2_8_zb;
  wire  [24:0] stage2_7_pr;
  wire  [24:0] stage2_7_sb;
  wire  [23:0] stage2_7_m0;
  wire  [23:0] stage2_7_m1;
  wire  [0:0] stage2_7_ms;
  wire  [23:0] stage2_7_mx;
  wire  [48:0] stage2_7_zl;
  wire  [0:0] stage2_7_zb;
  wire  [24:0] stage2_6_pr;
  wire  [24:0] stage2_6_sb;
  wire  [23:0] stage2_6_m0;
  wire  [23:0] stage2_6_m1;
  wire  [0:0] stage2_6_ms;
  wire  [23:0] stage2_6_mx;
  wire  [48:0] stage2_6_zl;
  wire  [0:0] stage2_6_zb;
  wire  [24:0] stage2_5_pr;
  wire  [24:0] stage2_5_sb;
  wire  [23:0] stage2_5_m0;
  wire  [23:0] stage2_5_m1;
  wire  [0:0] stage2_5_ms;
  wire  [23:0] stage2_5_mx;
  wire  [48:0] stage2_5_zl;
  wire  [0:0] stage2_5_zb;
  wire  [24:0] stage2_4_pr;
  wire  [24:0] stage2_4_sb;
  wire  [23:0] stage2_4_m0;
  wire  [23:0] stage2_4_m1;
  wire  [0:0] stage2_4_ms;
  wire  [23:0] stage2_4_mx;
  wire  [48:0] stage2_4_zl;
  wire  [0:0] stage2_4_zb;
  wire  [24:0] stage2_3_pr;
  wire  [24:0] stage2_3_sb;
  wire  [23:0] stage2_3_m0;
  wire  [23:0] stage2_3_m1;
  wire  [0:0] stage2_3_ms;
  wire  [23:0] stage2_3_mx;
  wire  [48:0] stage2_3_zl;
  wire  [0:0] stage2_3_zb;
  wire  [24:0] stage2_2_pr;
  wire  [24:0] stage2_2_sb;
  wire  [23:0] stage2_2_m0;
  wire  [23:0] stage2_2_m1;
  wire  [0:0] stage2_2_ms;
  wire  [23:0] stage2_2_mx;
  wire  [48:0] stage2_2_zl;
  wire  [0:0] stage2_2_zb;
  wire  [24:0] stage2_1_pr;
  wire  [24:0] stage2_1_sb;
  wire  [23:0] stage2_1_m0;
  wire  [23:0] stage2_1_m1;
  wire  [0:0] stage2_1_ms;
  wire  [23:0] stage2_1_mx;
  wire  [48:0] stage2_1_zl;
  wire  [0:0] stage2_1_zb;
  wire  [24:0] stage2_0_pr;
  wire  [24:0] stage2_0_sb;
  wire  [23:0] stage2_0_m0;
  wire  [23:0] stage2_0_m1;
  wire  [0:0] stage2_0_ms;
  wire  [23:0] stage2_0_mx;
  wire  [48:0] stage2_0_zl;
  wire  [0:0] stage2_0_zb;
  wire  [0:0] stage3_z_msb;
  wire  [24:0] anon_1008;
  wire  [26:0] anon_1009;
  wire  [25:0] anon_1010;
  wire  [26:0] anon_1011;
  wire  [0:0] anon_1012;
  wire  [23:0] stage4_fraction_data;
  wire  [0:0] stage4_s_least;
  wire  [0:0] stage4_s_guard;
  wire  [0:0] stage4_s_round;
  wire  [0:0] stage4_s_sticky;
  wire  [0:0] stage4_increment;
  wire  [0:0] anon_1026;
  wire  [0:0] anon_1027;
  wire  anon_1028;
  wire  [0:0] anon_1029;
  wire  stage5_exp_natural;
  wire  stage5_exp_underflow;
  wire  stage5_exp_overflow;
  wire  [7:0] stage5_exponent_in;
  wire  [22:0] stage5_fraction_in;
  wire  [7:0] stage5_exponent_i1;
  wire  [22:0] stage5_fraction_i1;
  wire  [7:0] stage5_exponent_di;
  wire  [22:0] stage5_fraction_di;
  wire  stage5_a_is_zero;
  wire  stage5_a_is_inf;
  wire  stage5_a_is_nan;
  wire  stage5_a_is_norm;
  wire  anon_1056;
  wire  anon_1057;
  wire  stage5_b_is_zero;
  wire  stage5_b_is_inf;
  wire  stage5_b_is_nan;
  wire  stage5_b_is_norm;
  wire  anon_1062;
  wire  anon_1063;
  wire  stage5_set_zero;
  wire  anon_1065;
  wire  anon_1066;
  wire  anon_1067;
  wire  anon_1068;
  wire  stage5_set_inf;
  wire  anon_1070;
  wire  anon_1071;
  wire  anon_1072;
  wire  anon_1073;
  wire  stage5_set_norm;
  wire  stage5_set_nan;
  wire  anon_1076;
  wire  anon_1077;
  wire  anon_1078;
  wire  anon_1079;
  wire  anon_1080;
  wire  anon_1081;
  wire  anon_1082;
  wire  anon_1083;
  wire  anon_1084;
  wire  [22:0] stage5_fraction_o0;
  wire  [7:0] stage5_exponent_o0;
  wire  [22:0] stage5_fraction_o1;
  wire  [7:0] stage5_exponent_o1;
  wire  [0:0] stage5_sign_o;
  wire  [22:0] stage5_fraction_o;
  wire  [7:0] stage5_exponent_o;
  wire  [31:0] stage5_result;
  // Resources
  // eq:11
  wire [7:0] eq_11_s0;
  assign eq_11_s0 = stage1_a_exponent_in;
  wire [7:0] eq_11_s1;
  assign eq_11_s1 = 8'd0;
  wire eq_11_d0;
  assign eq_11_d0 = eq_11_s0 == eq_11_s1;
  // eq:17
  wire [22:0] eq_17_s0;
  assign eq_17_s0 = stage1_a_fraction_in;
  wire [22:0] eq_17_s1;
  assign eq_17_s1 = 23'd0;
  wire eq_17_d0;
  assign eq_17_d0 = eq_17_s0 == eq_17_s1;
  // eq:21
  wire [7:0] eq_21_s0;
  assign eq_21_s0 = stage1_b_exponent_in;
  wire [7:0] eq_21_s1;
  assign eq_21_s1 = 8'd0;
  wire eq_21_d0;
  assign eq_21_d0 = eq_21_s0 == eq_21_s1;
  // eq:27
  wire [22:0] eq_27_s0;
  assign eq_27_s0 = stage1_b_fraction_in;
  wire [22:0] eq_27_s1;
  assign eq_27_s1 = 23'd0;
  wire eq_27_d0;
  assign eq_27_d0 = eq_27_s0 == eq_27_s1;
  // sub:29
  wire [9:0] sub_29_s0;
  assign sub_29_s0 = stage2_50_exponent_a_in;
  wire [7:0] sub_29_s1;
  assign sub_29_s1 = 8'd127;
  wire signed [9:0] sub_29_d0;
  assign sub_29_d0 = sub_29_s0 - sub_29_s1;
  // sub:31
  wire [9:0] sub_31_s0;
  assign sub_31_s0 = stage2_50_exponent_b_in;
  wire [7:0] sub_31_s1;
  assign sub_31_s1 = 8'd127;
  wire signed [9:0] sub_31_d0;
  assign sub_31_d0 = sub_31_s0 - sub_31_s1;
  // sub:34
  wire signed [9:0] sub_34_s0;
  assign sub_34_s0 = stage2_50_exponent_a_d;
  wire signed [9:0] sub_34_s1;
  assign sub_34_s1 = stage2_50_exponent_b_d;
  wire signed [9:0] sub_34_d0;
  assign sub_34_d0 = sub_34_s0 - sub_34_s1;
  // eq:37
  wire [7:0] eq_37_s0;
  assign eq_37_s0 = stage1_a_exponent;
  wire [7:0] eq_37_s1;
  assign eq_37_s1 = 8'd255;
  wire eq_37_d0;
  assign eq_37_d0 = eq_37_s0 == eq_37_s1;
  // eq:44
  wire [7:0] eq_44_s0;
  assign eq_44_s0 = stage1_b_exponent;
  wire [7:0] eq_44_s1;
  assign eq_44_s1 = 8'd255;
  wire eq_44_d0;
  assign eq_44_d0 = eq_44_s0 == eq_44_s1;
  // sub:51
  wire [24:0] sub_51_s0;
  assign sub_51_s0 = stage2_49_pr;
  wire [23:0] sub_51_s1;
  assign sub_51_s1 = stage2_di_50;
  wire [24:0] sub_51_d0;
  assign sub_51_d0 = sub_51_s0 - sub_51_s1;
  // sub:69
  wire [24:0] sub_69_s0;
  assign sub_69_s0 = stage2_48_pr;
  wire [23:0] sub_69_s1;
  assign sub_69_s1 = stage2_di_49;
  wire [24:0] sub_69_d0;
  assign sub_69_d0 = sub_69_s0 - sub_69_s1;
  // sub:87
  wire [24:0] sub_87_s0;
  assign sub_87_s0 = stage2_47_pr;
  wire [23:0] sub_87_s1;
  assign sub_87_s1 = stage2_di_48;
  wire [24:0] sub_87_d0;
  assign sub_87_d0 = sub_87_s0 - sub_87_s1;
  // sub:105
  wire [24:0] sub_105_s0;
  assign sub_105_s0 = stage2_46_pr;
  wire [23:0] sub_105_s1;
  assign sub_105_s1 = stage2_di_47;
  wire [24:0] sub_105_d0;
  assign sub_105_d0 = sub_105_s0 - sub_105_s1;
  // sub:123
  wire [24:0] sub_123_s0;
  assign sub_123_s0 = stage2_45_pr;
  wire [23:0] sub_123_s1;
  assign sub_123_s1 = stage2_di_46;
  wire [24:0] sub_123_d0;
  assign sub_123_d0 = sub_123_s0 - sub_123_s1;
  // sub:141
  wire [24:0] sub_141_s0;
  assign sub_141_s0 = stage2_44_pr;
  wire [23:0] sub_141_s1;
  assign sub_141_s1 = stage2_di_45;
  wire [24:0] sub_141_d0;
  assign sub_141_d0 = sub_141_s0 - sub_141_s1;
  // sub:159
  wire [24:0] sub_159_s0;
  assign sub_159_s0 = stage2_43_pr;
  wire [23:0] sub_159_s1;
  assign sub_159_s1 = stage2_di_44;
  wire [24:0] sub_159_d0;
  assign sub_159_d0 = sub_159_s0 - sub_159_s1;
  // sub:177
  wire [24:0] sub_177_s0;
  assign sub_177_s0 = stage2_42_pr;
  wire [23:0] sub_177_s1;
  assign sub_177_s1 = stage2_di_43;
  wire [24:0] sub_177_d0;
  assign sub_177_d0 = sub_177_s0 - sub_177_s1;
  // sub:195
  wire [24:0] sub_195_s0;
  assign sub_195_s0 = stage2_41_pr;
  wire [23:0] sub_195_s1;
  assign sub_195_s1 = stage2_di_42;
  wire [24:0] sub_195_d0;
  assign sub_195_d0 = sub_195_s0 - sub_195_s1;
  // sub:213
  wire [24:0] sub_213_s0;
  assign sub_213_s0 = stage2_40_pr;
  wire [23:0] sub_213_s1;
  assign sub_213_s1 = stage2_di_41;
  wire [24:0] sub_213_d0;
  assign sub_213_d0 = sub_213_s0 - sub_213_s1;
  // sub:231
  wire [24:0] sub_231_s0;
  assign sub_231_s0 = stage2_39_pr;
  wire [23:0] sub_231_s1;
  assign sub_231_s1 = stage2_di_40;
  wire [24:0] sub_231_d0;
  assign sub_231_d0 = sub_231_s0 - sub_231_s1;
  // sub:249
  wire [24:0] sub_249_s0;
  assign sub_249_s0 = stage2_38_pr;
  wire [23:0] sub_249_s1;
  assign sub_249_s1 = stage2_di_39;
  wire [24:0] sub_249_d0;
  assign sub_249_d0 = sub_249_s0 - sub_249_s1;
  // sub:267
  wire [24:0] sub_267_s0;
  assign sub_267_s0 = stage2_37_pr;
  wire [23:0] sub_267_s1;
  assign sub_267_s1 = stage2_di_38;
  wire [24:0] sub_267_d0;
  assign sub_267_d0 = sub_267_s0 - sub_267_s1;
  // sub:285
  wire [24:0] sub_285_s0;
  assign sub_285_s0 = stage2_36_pr;
  wire [23:0] sub_285_s1;
  assign sub_285_s1 = stage2_di_37;
  wire [24:0] sub_285_d0;
  assign sub_285_d0 = sub_285_s0 - sub_285_s1;
  // sub:303
  wire [24:0] sub_303_s0;
  assign sub_303_s0 = stage2_35_pr;
  wire [23:0] sub_303_s1;
  assign sub_303_s1 = stage2_di_36;
  wire [24:0] sub_303_d0;
  assign sub_303_d0 = sub_303_s0 - sub_303_s1;
  // sub:321
  wire [24:0] sub_321_s0;
  assign sub_321_s0 = stage2_34_pr;
  wire [23:0] sub_321_s1;
  assign sub_321_s1 = stage2_di_35;
  wire [24:0] sub_321_d0;
  assign sub_321_d0 = sub_321_s0 - sub_321_s1;
  // sub:339
  wire [24:0] sub_339_s0;
  assign sub_339_s0 = stage2_33_pr;
  wire [23:0] sub_339_s1;
  assign sub_339_s1 = stage2_di_34;
  wire [24:0] sub_339_d0;
  assign sub_339_d0 = sub_339_s0 - sub_339_s1;
  // sub:357
  wire [24:0] sub_357_s0;
  assign sub_357_s0 = stage2_32_pr;
  wire [23:0] sub_357_s1;
  assign sub_357_s1 = stage2_di_33;
  wire [24:0] sub_357_d0;
  assign sub_357_d0 = sub_357_s0 - sub_357_s1;
  // sub:375
  wire [24:0] sub_375_s0;
  assign sub_375_s0 = stage2_31_pr;
  wire [23:0] sub_375_s1;
  assign sub_375_s1 = stage2_di_32;
  wire [24:0] sub_375_d0;
  assign sub_375_d0 = sub_375_s0 - sub_375_s1;
  // sub:393
  wire [24:0] sub_393_s0;
  assign sub_393_s0 = stage2_30_pr;
  wire [23:0] sub_393_s1;
  assign sub_393_s1 = stage2_di_31;
  wire [24:0] sub_393_d0;
  assign sub_393_d0 = sub_393_s0 - sub_393_s1;
  // sub:411
  wire [24:0] sub_411_s0;
  assign sub_411_s0 = stage2_29_pr;
  wire [23:0] sub_411_s1;
  assign sub_411_s1 = stage2_di_30;
  wire [24:0] sub_411_d0;
  assign sub_411_d0 = sub_411_s0 - sub_411_s1;
  // sub:429
  wire [24:0] sub_429_s0;
  assign sub_429_s0 = stage2_28_pr;
  wire [23:0] sub_429_s1;
  assign sub_429_s1 = stage2_di_29;
  wire [24:0] sub_429_d0;
  assign sub_429_d0 = sub_429_s0 - sub_429_s1;
  // sub:447
  wire [24:0] sub_447_s0;
  assign sub_447_s0 = stage2_27_pr;
  wire [23:0] sub_447_s1;
  assign sub_447_s1 = stage2_di_28;
  wire [24:0] sub_447_d0;
  assign sub_447_d0 = sub_447_s0 - sub_447_s1;
  // sub:465
  wire [24:0] sub_465_s0;
  assign sub_465_s0 = stage2_26_pr;
  wire [23:0] sub_465_s1;
  assign sub_465_s1 = stage2_di_27;
  wire [24:0] sub_465_d0;
  assign sub_465_d0 = sub_465_s0 - sub_465_s1;
  // sub:483
  wire [24:0] sub_483_s0;
  assign sub_483_s0 = stage2_25_pr;
  wire [23:0] sub_483_s1;
  assign sub_483_s1 = stage2_di_26;
  wire [24:0] sub_483_d0;
  assign sub_483_d0 = sub_483_s0 - sub_483_s1;
  // sub:501
  wire [24:0] sub_501_s0;
  assign sub_501_s0 = stage2_24_pr;
  wire [23:0] sub_501_s1;
  assign sub_501_s1 = stage2_di_25;
  wire [24:0] sub_501_d0;
  assign sub_501_d0 = sub_501_s0 - sub_501_s1;
  // sub:519
  wire [24:0] sub_519_s0;
  assign sub_519_s0 = stage2_23_pr;
  wire [23:0] sub_519_s1;
  assign sub_519_s1 = stage2_di_24;
  wire [24:0] sub_519_d0;
  assign sub_519_d0 = sub_519_s0 - sub_519_s1;
  // sub:537
  wire [24:0] sub_537_s0;
  assign sub_537_s0 = stage2_22_pr;
  wire [23:0] sub_537_s1;
  assign sub_537_s1 = stage2_di_23;
  wire [24:0] sub_537_d0;
  assign sub_537_d0 = sub_537_s0 - sub_537_s1;
  // sub:555
  wire [24:0] sub_555_s0;
  assign sub_555_s0 = stage2_21_pr;
  wire [23:0] sub_555_s1;
  assign sub_555_s1 = stage2_di_22;
  wire [24:0] sub_555_d0;
  assign sub_555_d0 = sub_555_s0 - sub_555_s1;
  // sub:573
  wire [24:0] sub_573_s0;
  assign sub_573_s0 = stage2_20_pr;
  wire [23:0] sub_573_s1;
  assign sub_573_s1 = stage2_di_21;
  wire [24:0] sub_573_d0;
  assign sub_573_d0 = sub_573_s0 - sub_573_s1;
  // sub:591
  wire [24:0] sub_591_s0;
  assign sub_591_s0 = stage2_19_pr;
  wire [23:0] sub_591_s1;
  assign sub_591_s1 = stage2_di_20;
  wire [24:0] sub_591_d0;
  assign sub_591_d0 = sub_591_s0 - sub_591_s1;
  // sub:609
  wire [24:0] sub_609_s0;
  assign sub_609_s0 = stage2_18_pr;
  wire [23:0] sub_609_s1;
  assign sub_609_s1 = stage2_di_19;
  wire [24:0] sub_609_d0;
  assign sub_609_d0 = sub_609_s0 - sub_609_s1;
  // sub:627
  wire [24:0] sub_627_s0;
  assign sub_627_s0 = stage2_17_pr;
  wire [23:0] sub_627_s1;
  assign sub_627_s1 = stage2_di_18;
  wire [24:0] sub_627_d0;
  assign sub_627_d0 = sub_627_s0 - sub_627_s1;
  // sub:645
  wire [24:0] sub_645_s0;
  assign sub_645_s0 = stage2_16_pr;
  wire [23:0] sub_645_s1;
  assign sub_645_s1 = stage2_di_17;
  wire [24:0] sub_645_d0;
  assign sub_645_d0 = sub_645_s0 - sub_645_s1;
  // sub:663
  wire [24:0] sub_663_s0;
  assign sub_663_s0 = stage2_15_pr;
  wire [23:0] sub_663_s1;
  assign sub_663_s1 = stage2_di_16;
  wire [24:0] sub_663_d0;
  assign sub_663_d0 = sub_663_s0 - sub_663_s1;
  // sub:681
  wire [24:0] sub_681_s0;
  assign sub_681_s0 = stage2_14_pr;
  wire [23:0] sub_681_s1;
  assign sub_681_s1 = stage2_di_15;
  wire [24:0] sub_681_d0;
  assign sub_681_d0 = sub_681_s0 - sub_681_s1;
  // sub:699
  wire [24:0] sub_699_s0;
  assign sub_699_s0 = stage2_13_pr;
  wire [23:0] sub_699_s1;
  assign sub_699_s1 = stage2_di_14;
  wire [24:0] sub_699_d0;
  assign sub_699_d0 = sub_699_s0 - sub_699_s1;
  // sub:717
  wire [24:0] sub_717_s0;
  assign sub_717_s0 = stage2_12_pr;
  wire [23:0] sub_717_s1;
  assign sub_717_s1 = stage2_di_13;
  wire [24:0] sub_717_d0;
  assign sub_717_d0 = sub_717_s0 - sub_717_s1;
  // sub:735
  wire [24:0] sub_735_s0;
  assign sub_735_s0 = stage2_11_pr;
  wire [23:0] sub_735_s1;
  assign sub_735_s1 = stage2_di_12;
  wire [24:0] sub_735_d0;
  assign sub_735_d0 = sub_735_s0 - sub_735_s1;
  // sub:753
  wire [24:0] sub_753_s0;
  assign sub_753_s0 = stage2_10_pr;
  wire [23:0] sub_753_s1;
  assign sub_753_s1 = stage2_di_11;
  wire [24:0] sub_753_d0;
  assign sub_753_d0 = sub_753_s0 - sub_753_s1;
  // sub:771
  wire [24:0] sub_771_s0;
  assign sub_771_s0 = stage2_9_pr;
  wire [23:0] sub_771_s1;
  assign sub_771_s1 = stage2_di_10;
  wire [24:0] sub_771_d0;
  assign sub_771_d0 = sub_771_s0 - sub_771_s1;
  // sub:789
  wire [24:0] sub_789_s0;
  assign sub_789_s0 = stage2_8_pr;
  wire [23:0] sub_789_s1;
  assign sub_789_s1 = stage2_di_09;
  wire [24:0] sub_789_d0;
  assign sub_789_d0 = sub_789_s0 - sub_789_s1;
  // sub:807
  wire [24:0] sub_807_s0;
  assign sub_807_s0 = stage2_7_pr;
  wire [23:0] sub_807_s1;
  assign sub_807_s1 = stage2_di_08;
  wire [24:0] sub_807_d0;
  assign sub_807_d0 = sub_807_s0 - sub_807_s1;
  // sub:825
  wire [24:0] sub_825_s0;
  assign sub_825_s0 = stage2_6_pr;
  wire [23:0] sub_825_s1;
  assign sub_825_s1 = stage2_di_07;
  wire [24:0] sub_825_d0;
  assign sub_825_d0 = sub_825_s0 - sub_825_s1;
  // sub:843
  wire [24:0] sub_843_s0;
  assign sub_843_s0 = stage2_5_pr;
  wire [23:0] sub_843_s1;
  assign sub_843_s1 = stage2_di_06;
  wire [24:0] sub_843_d0;
  assign sub_843_d0 = sub_843_s0 - sub_843_s1;
  // sub:861
  wire [24:0] sub_861_s0;
  assign sub_861_s0 = stage2_4_pr;
  wire [23:0] sub_861_s1;
  assign sub_861_s1 = stage2_di_05;
  wire [24:0] sub_861_d0;
  assign sub_861_d0 = sub_861_s0 - sub_861_s1;
  // sub:879
  wire [24:0] sub_879_s0;
  assign sub_879_s0 = stage2_3_pr;
  wire [23:0] sub_879_s1;
  assign sub_879_s1 = stage2_di_04;
  wire [24:0] sub_879_d0;
  assign sub_879_d0 = sub_879_s0 - sub_879_s1;
  // sub:897
  wire [24:0] sub_897_s0;
  assign sub_897_s0 = stage2_2_pr;
  wire [23:0] sub_897_s1;
  assign sub_897_s1 = stage2_di_03;
  wire [24:0] sub_897_d0;
  assign sub_897_d0 = sub_897_s0 - sub_897_s1;
  // sub:915
  wire [24:0] sub_915_s0;
  assign sub_915_s0 = stage2_1_pr;
  wire [23:0] sub_915_s1;
  assign sub_915_s1 = stage2_di_02;
  wire [24:0] sub_915_d0;
  assign sub_915_d0 = sub_915_s0 - sub_915_s1;
  // sub:933
  wire [24:0] sub_933_s0;
  assign sub_933_s0 = stage2_0_pr;
  wire [23:0] sub_933_s1;
  assign sub_933_s1 = stage2_di_01;
  wire [24:0] sub_933_d0;
  assign sub_933_d0 = sub_933_s0 - sub_933_s1;
  // add:949
  wire signed [9:0] add_949_s0;
  assign add_949_s0 = stage2_exponent_01;
  wire [7:0] add_949_s1;
  assign add_949_s1 = 8'd127;
  wire signed [9:0] add_949_d0;
  assign add_949_d0 = add_949_s0 + add_949_s1;
  // sub:957
  wire signed [9:0] sub_957_s0;
  assign sub_957_s0 = stage2_exponent_00;
  wire [0:0] sub_957_s1;
  assign sub_957_s1 = anon_1012;
  wire signed [9:0] sub_957_d0;
  assign sub_957_d0 = sub_957_s0 - sub_957_s1;
  // add:973
  wire [23:0] add_973_s0;
  assign add_973_s0 = stage4_fraction_data;
  wire [0:0] add_973_s1;
  assign add_973_s1 = stage4_increment;
  wire [23:0] add_973_d0;
  assign add_973_d0 = add_973_s0 + add_973_s1;
  // eq:974
  wire [23:0] eq_974_s0;
  assign eq_974_s0 = stage4_fraction_data;
  wire [23:0] eq_974_s1;
  assign eq_974_s1 = 24'd16777215;
  wire eq_974_d0;
  assign eq_974_d0 = eq_974_s0 == eq_974_s1;
  // add:976
  wire signed [9:0] add_976_s0;
  assign add_976_s0 = stage3_exponent;
  wire [0:0] add_976_s1;
  assign add_976_s1 = anon_1029;
  wire signed [9:0] add_976_d0;
  assign add_976_d0 = add_976_s0 + add_976_s1;
  // gt:984
  wire signed [9:0] gt_984_s0;
  assign gt_984_s0 = stage4_exponent;
  wire signed [9:0] gt_984_s1;
  assign gt_984_s1 = 10'd0;
  wire gt_984_d0;
  assign gt_984_d0 = gt_984_s0 > gt_984_s1;
  // gte:986
  wire signed [9:0] gte_986_s0;
  assign gte_986_s0 = stage4_exponent;
  wire signed [9:0] gte_986_s1;
  assign gte_986_s1 = 10'd255;
  wire gte_986_d0;
  assign gte_986_d0 = gte_986_s0 >= gte_986_s1;
  // Insn wires
  wire  [0:0] insn_o_1_4_0;
  wire  [31:0] insn_o_1_5_0;
  wire  [7:0] insn_o_1_6_0;
  wire  [22:0] insn_o_1_7_0;
  wire  insn_o_1_8_0;
  wire  insn_o_1_9_0;
  wire  [0:0] insn_o_1_10_0;
  wire  [23:0] insn_o_1_11_0;
  wire  [7:0] insn_o_1_12_0;
  wire  insn_o_1_13_0;
  wire  insn_o_1_14_0;
  wire  insn_o_1_15_0;
  wire  [31:0] insn_o_1_16_0;
  wire  [7:0] insn_o_1_17_0;
  wire  [22:0] insn_o_1_18_0;
  wire  insn_o_1_19_0;
  wire  insn_o_1_20_0;
  wire  [0:0] insn_o_1_21_0;
  wire  [23:0] insn_o_1_22_0;
  wire  [7:0] insn_o_1_23_0;
  wire  insn_o_1_24_0;
  wire  insn_o_1_25_0;
  wire  insn_o_1_26_0;
  wire  [9:0] insn_o_1_28_0;
  wire  signed [9:0] insn_o_1_29_0;
  wire  [9:0] insn_o_1_30_0;
  wire  signed [9:0] insn_o_1_31_0;
  wire  [73:0] insn_o_1_32_0;
  wire  [23:0] insn_o_1_33_0;
  wire  signed [9:0] insn_o_1_34_0;
  wire  insn_o_1_35_0;
  wire  insn_o_1_36_0;
  wire  insn_o_1_37_0;
  wire  insn_o_1_38_0;
  wire  insn_o_1_39_0;
  wire  insn_o_1_40_0;
  wire  insn_o_1_41_0;
  wire  insn_o_1_42_0;
  wire  insn_o_1_43_0;
  wire  insn_o_1_44_0;
  wire  insn_o_1_45_0;
  wire  insn_o_1_46_0;
  wire  insn_o_1_47_0;
  wire  insn_o_1_48_0;
  wire  insn_o_1_49_0;
  wire  [24:0] insn_o_1_51_0;
  wire  [24:0] insn_o_1_52_0;
  wire  [23:0] insn_o_1_53_0;
  wire  [23:0] insn_o_1_54_0;
  wire  [0:0] insn_o_1_55_0;
  wire  [23:0] insn_o_1_56_0;
  wire  [48:0] insn_o_1_57_0;
  wire  [0:0] insn_o_1_58_0;
  wire  [73:0] insn_o_1_59_0;
  wire  [23:0] insn_o_1_60_0;
  wire  insn_o_1_61_0;
  wire  insn_o_1_62_0;
  wire  insn_o_1_63_0;
  wire  insn_o_1_64_0;
  wire  insn_o_1_65_0;
  wire  insn_o_1_66_0;
  wire  insn_o_1_67_0;
  wire  signed [9:0] insn_o_1_68_0;
  wire  [24:0] insn_o_1_70_0;
  wire  [24:0] insn_o_1_71_0;
  wire  [23:0] insn_o_1_72_0;
  wire  [23:0] insn_o_1_73_0;
  wire  [0:0] insn_o_1_74_0;
  wire  [23:0] insn_o_1_75_0;
  wire  [48:0] insn_o_1_76_0;
  wire  [0:0] insn_o_1_77_0;
  wire  [73:0] insn_o_1_78_0;
  wire  [23:0] insn_o_1_79_0;
  wire  insn_o_1_80_0;
  wire  insn_o_1_81_0;
  wire  insn_o_1_82_0;
  wire  insn_o_1_83_0;
  wire  insn_o_1_84_0;
  wire  insn_o_1_85_0;
  wire  insn_o_1_86_0;
  wire  signed [9:0] insn_o_1_87_0;
  wire  [24:0] insn_o_1_89_0;
  wire  [24:0] insn_o_1_90_0;
  wire  [23:0] insn_o_1_91_0;
  wire  [23:0] insn_o_1_92_0;
  wire  [0:0] insn_o_1_93_0;
  wire  [23:0] insn_o_1_94_0;
  wire  [48:0] insn_o_1_95_0;
  wire  [0:0] insn_o_1_96_0;
  wire  [73:0] insn_o_1_97_0;
  wire  [23:0] insn_o_1_98_0;
  wire  insn_o_1_99_0;
  wire  insn_o_1_100_0;
  wire  insn_o_1_101_0;
  wire  insn_o_1_102_0;
  wire  insn_o_1_103_0;
  wire  insn_o_1_104_0;
  wire  insn_o_1_105_0;
  wire  signed [9:0] insn_o_1_106_0;
  wire  [24:0] insn_o_1_108_0;
  wire  [24:0] insn_o_1_109_0;
  wire  [23:0] insn_o_1_110_0;
  wire  [23:0] insn_o_1_111_0;
  wire  [0:0] insn_o_1_112_0;
  wire  [23:0] insn_o_1_113_0;
  wire  [48:0] insn_o_1_114_0;
  wire  [0:0] insn_o_1_115_0;
  wire  [73:0] insn_o_1_116_0;
  wire  [23:0] insn_o_1_117_0;
  wire  insn_o_1_118_0;
  wire  insn_o_1_119_0;
  wire  insn_o_1_120_0;
  wire  insn_o_1_121_0;
  wire  insn_o_1_122_0;
  wire  insn_o_1_123_0;
  wire  insn_o_1_124_0;
  wire  signed [9:0] insn_o_1_125_0;
  wire  [24:0] insn_o_1_127_0;
  wire  [24:0] insn_o_1_128_0;
  wire  [23:0] insn_o_1_129_0;
  wire  [23:0] insn_o_1_130_0;
  wire  [0:0] insn_o_1_131_0;
  wire  [23:0] insn_o_1_132_0;
  wire  [48:0] insn_o_1_133_0;
  wire  [0:0] insn_o_1_134_0;
  wire  [73:0] insn_o_1_135_0;
  wire  [23:0] insn_o_1_136_0;
  wire  insn_o_1_137_0;
  wire  insn_o_1_138_0;
  wire  insn_o_1_139_0;
  wire  insn_o_1_140_0;
  wire  insn_o_1_141_0;
  wire  insn_o_1_142_0;
  wire  insn_o_1_143_0;
  wire  signed [9:0] insn_o_1_144_0;
  wire  [24:0] insn_o_1_146_0;
  wire  [24:0] insn_o_1_147_0;
  wire  [23:0] insn_o_1_148_0;
  wire  [23:0] insn_o_1_149_0;
  wire  [0:0] insn_o_1_150_0;
  wire  [23:0] insn_o_1_151_0;
  wire  [48:0] insn_o_1_152_0;
  wire  [0:0] insn_o_1_153_0;
  wire  [73:0] insn_o_1_154_0;
  wire  [23:0] insn_o_1_155_0;
  wire  insn_o_1_156_0;
  wire  insn_o_1_157_0;
  wire  insn_o_1_158_0;
  wire  insn_o_1_159_0;
  wire  insn_o_1_160_0;
  wire  insn_o_1_161_0;
  wire  insn_o_1_162_0;
  wire  signed [9:0] insn_o_1_163_0;
  wire  [24:0] insn_o_1_165_0;
  wire  [24:0] insn_o_1_166_0;
  wire  [23:0] insn_o_1_167_0;
  wire  [23:0] insn_o_1_168_0;
  wire  [0:0] insn_o_1_169_0;
  wire  [23:0] insn_o_1_170_0;
  wire  [48:0] insn_o_1_171_0;
  wire  [0:0] insn_o_1_172_0;
  wire  [73:0] insn_o_1_173_0;
  wire  [23:0] insn_o_1_174_0;
  wire  insn_o_1_175_0;
  wire  insn_o_1_176_0;
  wire  insn_o_1_177_0;
  wire  insn_o_1_178_0;
  wire  insn_o_1_179_0;
  wire  insn_o_1_180_0;
  wire  insn_o_1_181_0;
  wire  signed [9:0] insn_o_1_182_0;
  wire  [24:0] insn_o_1_184_0;
  wire  [24:0] insn_o_1_185_0;
  wire  [23:0] insn_o_1_186_0;
  wire  [23:0] insn_o_1_187_0;
  wire  [0:0] insn_o_1_188_0;
  wire  [23:0] insn_o_1_189_0;
  wire  [48:0] insn_o_1_190_0;
  wire  [0:0] insn_o_1_191_0;
  wire  [73:0] insn_o_1_192_0;
  wire  [23:0] insn_o_1_193_0;
  wire  insn_o_1_194_0;
  wire  insn_o_1_195_0;
  wire  insn_o_1_196_0;
  wire  insn_o_1_197_0;
  wire  insn_o_1_198_0;
  wire  insn_o_1_199_0;
  wire  insn_o_1_200_0;
  wire  signed [9:0] insn_o_1_201_0;
  wire  [24:0] insn_o_1_203_0;
  wire  [24:0] insn_o_1_204_0;
  wire  [23:0] insn_o_1_205_0;
  wire  [23:0] insn_o_1_206_0;
  wire  [0:0] insn_o_1_207_0;
  wire  [23:0] insn_o_1_208_0;
  wire  [48:0] insn_o_1_209_0;
  wire  [0:0] insn_o_1_210_0;
  wire  [73:0] insn_o_1_211_0;
  wire  [23:0] insn_o_1_212_0;
  wire  insn_o_1_213_0;
  wire  insn_o_1_214_0;
  wire  insn_o_1_215_0;
  wire  insn_o_1_216_0;
  wire  insn_o_1_217_0;
  wire  insn_o_1_218_0;
  wire  insn_o_1_219_0;
  wire  signed [9:0] insn_o_1_220_0;
  wire  [24:0] insn_o_1_222_0;
  wire  [24:0] insn_o_1_223_0;
  wire  [23:0] insn_o_1_224_0;
  wire  [23:0] insn_o_1_225_0;
  wire  [0:0] insn_o_1_226_0;
  wire  [23:0] insn_o_1_227_0;
  wire  [48:0] insn_o_1_228_0;
  wire  [0:0] insn_o_1_229_0;
  wire  [73:0] insn_o_1_230_0;
  wire  [23:0] insn_o_1_231_0;
  wire  insn_o_1_232_0;
  wire  insn_o_1_233_0;
  wire  insn_o_1_234_0;
  wire  insn_o_1_235_0;
  wire  insn_o_1_236_0;
  wire  insn_o_1_237_0;
  wire  insn_o_1_238_0;
  wire  signed [9:0] insn_o_1_239_0;
  wire  [24:0] insn_o_1_241_0;
  wire  [24:0] insn_o_1_242_0;
  wire  [23:0] insn_o_1_243_0;
  wire  [23:0] insn_o_1_244_0;
  wire  [0:0] insn_o_1_245_0;
  wire  [23:0] insn_o_1_246_0;
  wire  [48:0] insn_o_1_247_0;
  wire  [0:0] insn_o_1_248_0;
  wire  [73:0] insn_o_1_249_0;
  wire  [23:0] insn_o_1_250_0;
  wire  insn_o_1_251_0;
  wire  insn_o_1_252_0;
  wire  insn_o_1_253_0;
  wire  insn_o_1_254_0;
  wire  insn_o_1_255_0;
  wire  insn_o_1_256_0;
  wire  insn_o_1_257_0;
  wire  signed [9:0] insn_o_1_258_0;
  wire  [24:0] insn_o_1_260_0;
  wire  [24:0] insn_o_1_261_0;
  wire  [23:0] insn_o_1_262_0;
  wire  [23:0] insn_o_1_263_0;
  wire  [0:0] insn_o_1_264_0;
  wire  [23:0] insn_o_1_265_0;
  wire  [48:0] insn_o_1_266_0;
  wire  [0:0] insn_o_1_267_0;
  wire  [73:0] insn_o_1_268_0;
  wire  [23:0] insn_o_1_269_0;
  wire  insn_o_1_270_0;
  wire  insn_o_1_271_0;
  wire  insn_o_1_272_0;
  wire  insn_o_1_273_0;
  wire  insn_o_1_274_0;
  wire  insn_o_1_275_0;
  wire  insn_o_1_276_0;
  wire  signed [9:0] insn_o_1_277_0;
  wire  [24:0] insn_o_1_279_0;
  wire  [24:0] insn_o_1_280_0;
  wire  [23:0] insn_o_1_281_0;
  wire  [23:0] insn_o_1_282_0;
  wire  [0:0] insn_o_1_283_0;
  wire  [23:0] insn_o_1_284_0;
  wire  [48:0] insn_o_1_285_0;
  wire  [0:0] insn_o_1_286_0;
  wire  [73:0] insn_o_1_287_0;
  wire  [23:0] insn_o_1_288_0;
  wire  insn_o_1_289_0;
  wire  insn_o_1_290_0;
  wire  insn_o_1_291_0;
  wire  insn_o_1_292_0;
  wire  insn_o_1_293_0;
  wire  insn_o_1_294_0;
  wire  insn_o_1_295_0;
  wire  signed [9:0] insn_o_1_296_0;
  wire  [24:0] insn_o_1_298_0;
  wire  [24:0] insn_o_1_299_0;
  wire  [23:0] insn_o_1_300_0;
  wire  [23:0] insn_o_1_301_0;
  wire  [0:0] insn_o_1_302_0;
  wire  [23:0] insn_o_1_303_0;
  wire  [48:0] insn_o_1_304_0;
  wire  [0:0] insn_o_1_305_0;
  wire  [73:0] insn_o_1_306_0;
  wire  [23:0] insn_o_1_307_0;
  wire  insn_o_1_308_0;
  wire  insn_o_1_309_0;
  wire  insn_o_1_310_0;
  wire  insn_o_1_311_0;
  wire  insn_o_1_312_0;
  wire  insn_o_1_313_0;
  wire  insn_o_1_314_0;
  wire  signed [9:0] insn_o_1_315_0;
  wire  [24:0] insn_o_1_317_0;
  wire  [24:0] insn_o_1_318_0;
  wire  [23:0] insn_o_1_319_0;
  wire  [23:0] insn_o_1_320_0;
  wire  [0:0] insn_o_1_321_0;
  wire  [23:0] insn_o_1_322_0;
  wire  [48:0] insn_o_1_323_0;
  wire  [0:0] insn_o_1_324_0;
  wire  [73:0] insn_o_1_325_0;
  wire  [23:0] insn_o_1_326_0;
  wire  insn_o_1_327_0;
  wire  insn_o_1_328_0;
  wire  insn_o_1_329_0;
  wire  insn_o_1_330_0;
  wire  insn_o_1_331_0;
  wire  insn_o_1_332_0;
  wire  insn_o_1_333_0;
  wire  signed [9:0] insn_o_1_334_0;
  wire  [24:0] insn_o_1_336_0;
  wire  [24:0] insn_o_1_337_0;
  wire  [23:0] insn_o_1_338_0;
  wire  [23:0] insn_o_1_339_0;
  wire  [0:0] insn_o_1_340_0;
  wire  [23:0] insn_o_1_341_0;
  wire  [48:0] insn_o_1_342_0;
  wire  [0:0] insn_o_1_343_0;
  wire  [73:0] insn_o_1_344_0;
  wire  [23:0] insn_o_1_345_0;
  wire  insn_o_1_346_0;
  wire  insn_o_1_347_0;
  wire  insn_o_1_348_0;
  wire  insn_o_1_349_0;
  wire  insn_o_1_350_0;
  wire  insn_o_1_351_0;
  wire  insn_o_1_352_0;
  wire  signed [9:0] insn_o_1_353_0;
  wire  [24:0] insn_o_1_355_0;
  wire  [24:0] insn_o_1_356_0;
  wire  [23:0] insn_o_1_357_0;
  wire  [23:0] insn_o_1_358_0;
  wire  [0:0] insn_o_1_359_0;
  wire  [23:0] insn_o_1_360_0;
  wire  [48:0] insn_o_1_361_0;
  wire  [0:0] insn_o_1_362_0;
  wire  [73:0] insn_o_1_363_0;
  wire  [23:0] insn_o_1_364_0;
  wire  insn_o_1_365_0;
  wire  insn_o_1_366_0;
  wire  insn_o_1_367_0;
  wire  insn_o_1_368_0;
  wire  insn_o_1_369_0;
  wire  insn_o_1_370_0;
  wire  insn_o_1_371_0;
  wire  signed [9:0] insn_o_1_372_0;
  wire  [24:0] insn_o_1_374_0;
  wire  [24:0] insn_o_1_375_0;
  wire  [23:0] insn_o_1_376_0;
  wire  [23:0] insn_o_1_377_0;
  wire  [0:0] insn_o_1_378_0;
  wire  [23:0] insn_o_1_379_0;
  wire  [48:0] insn_o_1_380_0;
  wire  [0:0] insn_o_1_381_0;
  wire  [73:0] insn_o_1_382_0;
  wire  [23:0] insn_o_1_383_0;
  wire  insn_o_1_384_0;
  wire  insn_o_1_385_0;
  wire  insn_o_1_386_0;
  wire  insn_o_1_387_0;
  wire  insn_o_1_388_0;
  wire  insn_o_1_389_0;
  wire  insn_o_1_390_0;
  wire  signed [9:0] insn_o_1_391_0;
  wire  [24:0] insn_o_1_393_0;
  wire  [24:0] insn_o_1_394_0;
  wire  [23:0] insn_o_1_395_0;
  wire  [23:0] insn_o_1_396_0;
  wire  [0:0] insn_o_1_397_0;
  wire  [23:0] insn_o_1_398_0;
  wire  [48:0] insn_o_1_399_0;
  wire  [0:0] insn_o_1_400_0;
  wire  [73:0] insn_o_1_401_0;
  wire  [23:0] insn_o_1_402_0;
  wire  insn_o_1_403_0;
  wire  insn_o_1_404_0;
  wire  insn_o_1_405_0;
  wire  insn_o_1_406_0;
  wire  insn_o_1_407_0;
  wire  insn_o_1_408_0;
  wire  insn_o_1_409_0;
  wire  signed [9:0] insn_o_1_410_0;
  wire  [24:0] insn_o_1_412_0;
  wire  [24:0] insn_o_1_413_0;
  wire  [23:0] insn_o_1_414_0;
  wire  [23:0] insn_o_1_415_0;
  wire  [0:0] insn_o_1_416_0;
  wire  [23:0] insn_o_1_417_0;
  wire  [48:0] insn_o_1_418_0;
  wire  [0:0] insn_o_1_419_0;
  wire  [73:0] insn_o_1_420_0;
  wire  [23:0] insn_o_1_421_0;
  wire  insn_o_1_422_0;
  wire  insn_o_1_423_0;
  wire  insn_o_1_424_0;
  wire  insn_o_1_425_0;
  wire  insn_o_1_426_0;
  wire  insn_o_1_427_0;
  wire  insn_o_1_428_0;
  wire  signed [9:0] insn_o_1_429_0;
  wire  [24:0] insn_o_1_431_0;
  wire  [24:0] insn_o_1_432_0;
  wire  [23:0] insn_o_1_433_0;
  wire  [23:0] insn_o_1_434_0;
  wire  [0:0] insn_o_1_435_0;
  wire  [23:0] insn_o_1_436_0;
  wire  [48:0] insn_o_1_437_0;
  wire  [0:0] insn_o_1_438_0;
  wire  [73:0] insn_o_1_439_0;
  wire  [23:0] insn_o_1_440_0;
  wire  insn_o_1_441_0;
  wire  insn_o_1_442_0;
  wire  insn_o_1_443_0;
  wire  insn_o_1_444_0;
  wire  insn_o_1_445_0;
  wire  insn_o_1_446_0;
  wire  insn_o_1_447_0;
  wire  signed [9:0] insn_o_1_448_0;
  wire  [24:0] insn_o_1_450_0;
  wire  [24:0] insn_o_1_451_0;
  wire  [23:0] insn_o_1_452_0;
  wire  [23:0] insn_o_1_453_0;
  wire  [0:0] insn_o_1_454_0;
  wire  [23:0] insn_o_1_455_0;
  wire  [48:0] insn_o_1_456_0;
  wire  [0:0] insn_o_1_457_0;
  wire  [73:0] insn_o_1_458_0;
  wire  [23:0] insn_o_1_459_0;
  wire  insn_o_1_460_0;
  wire  insn_o_1_461_0;
  wire  insn_o_1_462_0;
  wire  insn_o_1_463_0;
  wire  insn_o_1_464_0;
  wire  insn_o_1_465_0;
  wire  insn_o_1_466_0;
  wire  signed [9:0] insn_o_1_467_0;
  wire  [24:0] insn_o_1_469_0;
  wire  [24:0] insn_o_1_470_0;
  wire  [23:0] insn_o_1_471_0;
  wire  [23:0] insn_o_1_472_0;
  wire  [0:0] insn_o_1_473_0;
  wire  [23:0] insn_o_1_474_0;
  wire  [48:0] insn_o_1_475_0;
  wire  [0:0] insn_o_1_476_0;
  wire  [73:0] insn_o_1_477_0;
  wire  [23:0] insn_o_1_478_0;
  wire  insn_o_1_479_0;
  wire  insn_o_1_480_0;
  wire  insn_o_1_481_0;
  wire  insn_o_1_482_0;
  wire  insn_o_1_483_0;
  wire  insn_o_1_484_0;
  wire  insn_o_1_485_0;
  wire  signed [9:0] insn_o_1_486_0;
  wire  [24:0] insn_o_1_488_0;
  wire  [24:0] insn_o_1_489_0;
  wire  [23:0] insn_o_1_490_0;
  wire  [23:0] insn_o_1_491_0;
  wire  [0:0] insn_o_1_492_0;
  wire  [23:0] insn_o_1_493_0;
  wire  [48:0] insn_o_1_494_0;
  wire  [0:0] insn_o_1_495_0;
  wire  [73:0] insn_o_1_496_0;
  wire  [23:0] insn_o_1_497_0;
  wire  insn_o_1_498_0;
  wire  insn_o_1_499_0;
  wire  insn_o_1_500_0;
  wire  insn_o_1_501_0;
  wire  insn_o_1_502_0;
  wire  insn_o_1_503_0;
  wire  insn_o_1_504_0;
  wire  signed [9:0] insn_o_1_505_0;
  wire  [24:0] insn_o_1_507_0;
  wire  [24:0] insn_o_1_508_0;
  wire  [23:0] insn_o_1_509_0;
  wire  [23:0] insn_o_1_510_0;
  wire  [0:0] insn_o_1_511_0;
  wire  [23:0] insn_o_1_512_0;
  wire  [48:0] insn_o_1_513_0;
  wire  [0:0] insn_o_1_514_0;
  wire  [73:0] insn_o_1_515_0;
  wire  [23:0] insn_o_1_516_0;
  wire  insn_o_1_517_0;
  wire  insn_o_1_518_0;
  wire  insn_o_1_519_0;
  wire  insn_o_1_520_0;
  wire  insn_o_1_521_0;
  wire  insn_o_1_522_0;
  wire  insn_o_1_523_0;
  wire  signed [9:0] insn_o_1_524_0;
  wire  [24:0] insn_o_1_526_0;
  wire  [24:0] insn_o_1_527_0;
  wire  [23:0] insn_o_1_528_0;
  wire  [23:0] insn_o_1_529_0;
  wire  [0:0] insn_o_1_530_0;
  wire  [23:0] insn_o_1_531_0;
  wire  [48:0] insn_o_1_532_0;
  wire  [0:0] insn_o_1_533_0;
  wire  [73:0] insn_o_1_534_0;
  wire  [23:0] insn_o_1_535_0;
  wire  insn_o_1_536_0;
  wire  insn_o_1_537_0;
  wire  insn_o_1_538_0;
  wire  insn_o_1_539_0;
  wire  insn_o_1_540_0;
  wire  insn_o_1_541_0;
  wire  insn_o_1_542_0;
  wire  signed [9:0] insn_o_1_543_0;
  wire  [24:0] insn_o_1_545_0;
  wire  [24:0] insn_o_1_546_0;
  wire  [23:0] insn_o_1_547_0;
  wire  [23:0] insn_o_1_548_0;
  wire  [0:0] insn_o_1_549_0;
  wire  [23:0] insn_o_1_550_0;
  wire  [48:0] insn_o_1_551_0;
  wire  [0:0] insn_o_1_552_0;
  wire  [73:0] insn_o_1_553_0;
  wire  [23:0] insn_o_1_554_0;
  wire  insn_o_1_555_0;
  wire  insn_o_1_556_0;
  wire  insn_o_1_557_0;
  wire  insn_o_1_558_0;
  wire  insn_o_1_559_0;
  wire  insn_o_1_560_0;
  wire  insn_o_1_561_0;
  wire  signed [9:0] insn_o_1_562_0;
  wire  [24:0] insn_o_1_564_0;
  wire  [24:0] insn_o_1_565_0;
  wire  [23:0] insn_o_1_566_0;
  wire  [23:0] insn_o_1_567_0;
  wire  [0:0] insn_o_1_568_0;
  wire  [23:0] insn_o_1_569_0;
  wire  [48:0] insn_o_1_570_0;
  wire  [0:0] insn_o_1_571_0;
  wire  [73:0] insn_o_1_572_0;
  wire  [23:0] insn_o_1_573_0;
  wire  insn_o_1_574_0;
  wire  insn_o_1_575_0;
  wire  insn_o_1_576_0;
  wire  insn_o_1_577_0;
  wire  insn_o_1_578_0;
  wire  insn_o_1_579_0;
  wire  insn_o_1_580_0;
  wire  signed [9:0] insn_o_1_581_0;
  wire  [24:0] insn_o_1_583_0;
  wire  [24:0] insn_o_1_584_0;
  wire  [23:0] insn_o_1_585_0;
  wire  [23:0] insn_o_1_586_0;
  wire  [0:0] insn_o_1_587_0;
  wire  [23:0] insn_o_1_588_0;
  wire  [48:0] insn_o_1_589_0;
  wire  [0:0] insn_o_1_590_0;
  wire  [73:0] insn_o_1_591_0;
  wire  [23:0] insn_o_1_592_0;
  wire  insn_o_1_593_0;
  wire  insn_o_1_594_0;
  wire  insn_o_1_595_0;
  wire  insn_o_1_596_0;
  wire  insn_o_1_597_0;
  wire  insn_o_1_598_0;
  wire  insn_o_1_599_0;
  wire  signed [9:0] insn_o_1_600_0;
  wire  [24:0] insn_o_1_602_0;
  wire  [24:0] insn_o_1_603_0;
  wire  [23:0] insn_o_1_604_0;
  wire  [23:0] insn_o_1_605_0;
  wire  [0:0] insn_o_1_606_0;
  wire  [23:0] insn_o_1_607_0;
  wire  [48:0] insn_o_1_608_0;
  wire  [0:0] insn_o_1_609_0;
  wire  [73:0] insn_o_1_610_0;
  wire  [23:0] insn_o_1_611_0;
  wire  insn_o_1_612_0;
  wire  insn_o_1_613_0;
  wire  insn_o_1_614_0;
  wire  insn_o_1_615_0;
  wire  insn_o_1_616_0;
  wire  insn_o_1_617_0;
  wire  insn_o_1_618_0;
  wire  signed [9:0] insn_o_1_619_0;
  wire  [24:0] insn_o_1_621_0;
  wire  [24:0] insn_o_1_622_0;
  wire  [23:0] insn_o_1_623_0;
  wire  [23:0] insn_o_1_624_0;
  wire  [0:0] insn_o_1_625_0;
  wire  [23:0] insn_o_1_626_0;
  wire  [48:0] insn_o_1_627_0;
  wire  [0:0] insn_o_1_628_0;
  wire  [73:0] insn_o_1_629_0;
  wire  [23:0] insn_o_1_630_0;
  wire  insn_o_1_631_0;
  wire  insn_o_1_632_0;
  wire  insn_o_1_633_0;
  wire  insn_o_1_634_0;
  wire  insn_o_1_635_0;
  wire  insn_o_1_636_0;
  wire  insn_o_1_637_0;
  wire  signed [9:0] insn_o_1_638_0;
  wire  [24:0] insn_o_1_640_0;
  wire  [24:0] insn_o_1_641_0;
  wire  [23:0] insn_o_1_642_0;
  wire  [23:0] insn_o_1_643_0;
  wire  [0:0] insn_o_1_644_0;
  wire  [23:0] insn_o_1_645_0;
  wire  [48:0] insn_o_1_646_0;
  wire  [0:0] insn_o_1_647_0;
  wire  [73:0] insn_o_1_648_0;
  wire  [23:0] insn_o_1_649_0;
  wire  insn_o_1_650_0;
  wire  insn_o_1_651_0;
  wire  insn_o_1_652_0;
  wire  insn_o_1_653_0;
  wire  insn_o_1_654_0;
  wire  insn_o_1_655_0;
  wire  insn_o_1_656_0;
  wire  signed [9:0] insn_o_1_657_0;
  wire  [24:0] insn_o_1_659_0;
  wire  [24:0] insn_o_1_660_0;
  wire  [23:0] insn_o_1_661_0;
  wire  [23:0] insn_o_1_662_0;
  wire  [0:0] insn_o_1_663_0;
  wire  [23:0] insn_o_1_664_0;
  wire  [48:0] insn_o_1_665_0;
  wire  [0:0] insn_o_1_666_0;
  wire  [73:0] insn_o_1_667_0;
  wire  [23:0] insn_o_1_668_0;
  wire  insn_o_1_669_0;
  wire  insn_o_1_670_0;
  wire  insn_o_1_671_0;
  wire  insn_o_1_672_0;
  wire  insn_o_1_673_0;
  wire  insn_o_1_674_0;
  wire  insn_o_1_675_0;
  wire  signed [9:0] insn_o_1_676_0;
  wire  [24:0] insn_o_1_678_0;
  wire  [24:0] insn_o_1_679_0;
  wire  [23:0] insn_o_1_680_0;
  wire  [23:0] insn_o_1_681_0;
  wire  [0:0] insn_o_1_682_0;
  wire  [23:0] insn_o_1_683_0;
  wire  [48:0] insn_o_1_684_0;
  wire  [0:0] insn_o_1_685_0;
  wire  [73:0] insn_o_1_686_0;
  wire  [23:0] insn_o_1_687_0;
  wire  insn_o_1_688_0;
  wire  insn_o_1_689_0;
  wire  insn_o_1_690_0;
  wire  insn_o_1_691_0;
  wire  insn_o_1_692_0;
  wire  insn_o_1_693_0;
  wire  insn_o_1_694_0;
  wire  signed [9:0] insn_o_1_695_0;
  wire  [24:0] insn_o_1_697_0;
  wire  [24:0] insn_o_1_698_0;
  wire  [23:0] insn_o_1_699_0;
  wire  [23:0] insn_o_1_700_0;
  wire  [0:0] insn_o_1_701_0;
  wire  [23:0] insn_o_1_702_0;
  wire  [48:0] insn_o_1_703_0;
  wire  [0:0] insn_o_1_704_0;
  wire  [73:0] insn_o_1_705_0;
  wire  [23:0] insn_o_1_706_0;
  wire  insn_o_1_707_0;
  wire  insn_o_1_708_0;
  wire  insn_o_1_709_0;
  wire  insn_o_1_710_0;
  wire  insn_o_1_711_0;
  wire  insn_o_1_712_0;
  wire  insn_o_1_713_0;
  wire  signed [9:0] insn_o_1_714_0;
  wire  [24:0] insn_o_1_716_0;
  wire  [24:0] insn_o_1_717_0;
  wire  [23:0] insn_o_1_718_0;
  wire  [23:0] insn_o_1_719_0;
  wire  [0:0] insn_o_1_720_0;
  wire  [23:0] insn_o_1_721_0;
  wire  [48:0] insn_o_1_722_0;
  wire  [0:0] insn_o_1_723_0;
  wire  [73:0] insn_o_1_724_0;
  wire  [23:0] insn_o_1_725_0;
  wire  insn_o_1_726_0;
  wire  insn_o_1_727_0;
  wire  insn_o_1_728_0;
  wire  insn_o_1_729_0;
  wire  insn_o_1_730_0;
  wire  insn_o_1_731_0;
  wire  insn_o_1_732_0;
  wire  signed [9:0] insn_o_1_733_0;
  wire  [24:0] insn_o_1_735_0;
  wire  [24:0] insn_o_1_736_0;
  wire  [23:0] insn_o_1_737_0;
  wire  [23:0] insn_o_1_738_0;
  wire  [0:0] insn_o_1_739_0;
  wire  [23:0] insn_o_1_740_0;
  wire  [48:0] insn_o_1_741_0;
  wire  [0:0] insn_o_1_742_0;
  wire  [73:0] insn_o_1_743_0;
  wire  [23:0] insn_o_1_744_0;
  wire  insn_o_1_745_0;
  wire  insn_o_1_746_0;
  wire  insn_o_1_747_0;
  wire  insn_o_1_748_0;
  wire  insn_o_1_749_0;
  wire  insn_o_1_750_0;
  wire  insn_o_1_751_0;
  wire  signed [9:0] insn_o_1_752_0;
  wire  [24:0] insn_o_1_754_0;
  wire  [24:0] insn_o_1_755_0;
  wire  [23:0] insn_o_1_756_0;
  wire  [23:0] insn_o_1_757_0;
  wire  [0:0] insn_o_1_758_0;
  wire  [23:0] insn_o_1_759_0;
  wire  [48:0] insn_o_1_760_0;
  wire  [0:0] insn_o_1_761_0;
  wire  [73:0] insn_o_1_762_0;
  wire  [23:0] insn_o_1_763_0;
  wire  insn_o_1_764_0;
  wire  insn_o_1_765_0;
  wire  insn_o_1_766_0;
  wire  insn_o_1_767_0;
  wire  insn_o_1_768_0;
  wire  insn_o_1_769_0;
  wire  insn_o_1_770_0;
  wire  signed [9:0] insn_o_1_771_0;
  wire  [24:0] insn_o_1_773_0;
  wire  [24:0] insn_o_1_774_0;
  wire  [23:0] insn_o_1_775_0;
  wire  [23:0] insn_o_1_776_0;
  wire  [0:0] insn_o_1_777_0;
  wire  [23:0] insn_o_1_778_0;
  wire  [48:0] insn_o_1_779_0;
  wire  [0:0] insn_o_1_780_0;
  wire  [73:0] insn_o_1_781_0;
  wire  [23:0] insn_o_1_782_0;
  wire  insn_o_1_783_0;
  wire  insn_o_1_784_0;
  wire  insn_o_1_785_0;
  wire  insn_o_1_786_0;
  wire  insn_o_1_787_0;
  wire  insn_o_1_788_0;
  wire  insn_o_1_789_0;
  wire  signed [9:0] insn_o_1_790_0;
  wire  [24:0] insn_o_1_792_0;
  wire  [24:0] insn_o_1_793_0;
  wire  [23:0] insn_o_1_794_0;
  wire  [23:0] insn_o_1_795_0;
  wire  [0:0] insn_o_1_796_0;
  wire  [23:0] insn_o_1_797_0;
  wire  [48:0] insn_o_1_798_0;
  wire  [0:0] insn_o_1_799_0;
  wire  [73:0] insn_o_1_800_0;
  wire  [23:0] insn_o_1_801_0;
  wire  insn_o_1_802_0;
  wire  insn_o_1_803_0;
  wire  insn_o_1_804_0;
  wire  insn_o_1_805_0;
  wire  insn_o_1_806_0;
  wire  insn_o_1_807_0;
  wire  insn_o_1_808_0;
  wire  signed [9:0] insn_o_1_809_0;
  wire  [24:0] insn_o_1_811_0;
  wire  [24:0] insn_o_1_812_0;
  wire  [23:0] insn_o_1_813_0;
  wire  [23:0] insn_o_1_814_0;
  wire  [0:0] insn_o_1_815_0;
  wire  [23:0] insn_o_1_816_0;
  wire  [48:0] insn_o_1_817_0;
  wire  [0:0] insn_o_1_818_0;
  wire  [73:0] insn_o_1_819_0;
  wire  [23:0] insn_o_1_820_0;
  wire  insn_o_1_821_0;
  wire  insn_o_1_822_0;
  wire  insn_o_1_823_0;
  wire  insn_o_1_824_0;
  wire  insn_o_1_825_0;
  wire  insn_o_1_826_0;
  wire  insn_o_1_827_0;
  wire  signed [9:0] insn_o_1_828_0;
  wire  [24:0] insn_o_1_830_0;
  wire  [24:0] insn_o_1_831_0;
  wire  [23:0] insn_o_1_832_0;
  wire  [23:0] insn_o_1_833_0;
  wire  [0:0] insn_o_1_834_0;
  wire  [23:0] insn_o_1_835_0;
  wire  [48:0] insn_o_1_836_0;
  wire  [0:0] insn_o_1_837_0;
  wire  [73:0] insn_o_1_838_0;
  wire  [23:0] insn_o_1_839_0;
  wire  insn_o_1_840_0;
  wire  insn_o_1_841_0;
  wire  insn_o_1_842_0;
  wire  insn_o_1_843_0;
  wire  insn_o_1_844_0;
  wire  insn_o_1_845_0;
  wire  insn_o_1_846_0;
  wire  signed [9:0] insn_o_1_847_0;
  wire  [24:0] insn_o_1_849_0;
  wire  [24:0] insn_o_1_850_0;
  wire  [23:0] insn_o_1_851_0;
  wire  [23:0] insn_o_1_852_0;
  wire  [0:0] insn_o_1_853_0;
  wire  [23:0] insn_o_1_854_0;
  wire  [48:0] insn_o_1_855_0;
  wire  [0:0] insn_o_1_856_0;
  wire  [73:0] insn_o_1_857_0;
  wire  [23:0] insn_o_1_858_0;
  wire  insn_o_1_859_0;
  wire  insn_o_1_860_0;
  wire  insn_o_1_861_0;
  wire  insn_o_1_862_0;
  wire  insn_o_1_863_0;
  wire  insn_o_1_864_0;
  wire  insn_o_1_865_0;
  wire  signed [9:0] insn_o_1_866_0;
  wire  [24:0] insn_o_1_868_0;
  wire  [24:0] insn_o_1_869_0;
  wire  [23:0] insn_o_1_870_0;
  wire  [23:0] insn_o_1_871_0;
  wire  [0:0] insn_o_1_872_0;
  wire  [23:0] insn_o_1_873_0;
  wire  [48:0] insn_o_1_874_0;
  wire  [0:0] insn_o_1_875_0;
  wire  [73:0] insn_o_1_876_0;
  wire  [23:0] insn_o_1_877_0;
  wire  insn_o_1_878_0;
  wire  insn_o_1_879_0;
  wire  insn_o_1_880_0;
  wire  insn_o_1_881_0;
  wire  insn_o_1_882_0;
  wire  insn_o_1_883_0;
  wire  insn_o_1_884_0;
  wire  signed [9:0] insn_o_1_885_0;
  wire  [24:0] insn_o_1_887_0;
  wire  [24:0] insn_o_1_888_0;
  wire  [23:0] insn_o_1_889_0;
  wire  [23:0] insn_o_1_890_0;
  wire  [0:0] insn_o_1_891_0;
  wire  [23:0] insn_o_1_892_0;
  wire  [48:0] insn_o_1_893_0;
  wire  [0:0] insn_o_1_894_0;
  wire  [73:0] insn_o_1_895_0;
  wire  [23:0] insn_o_1_896_0;
  wire  insn_o_1_897_0;
  wire  insn_o_1_898_0;
  wire  insn_o_1_899_0;
  wire  insn_o_1_900_0;
  wire  insn_o_1_901_0;
  wire  insn_o_1_902_0;
  wire  insn_o_1_903_0;
  wire  signed [9:0] insn_o_1_904_0;
  wire  [24:0] insn_o_1_906_0;
  wire  [24:0] insn_o_1_907_0;
  wire  [23:0] insn_o_1_908_0;
  wire  [23:0] insn_o_1_909_0;
  wire  [0:0] insn_o_1_910_0;
  wire  [23:0] insn_o_1_911_0;
  wire  [48:0] insn_o_1_912_0;
  wire  [0:0] insn_o_1_913_0;
  wire  [73:0] insn_o_1_914_0;
  wire  [23:0] insn_o_1_915_0;
  wire  insn_o_1_916_0;
  wire  insn_o_1_917_0;
  wire  insn_o_1_918_0;
  wire  insn_o_1_919_0;
  wire  insn_o_1_920_0;
  wire  insn_o_1_921_0;
  wire  insn_o_1_922_0;
  wire  signed [9:0] insn_o_1_923_0;
  wire  [24:0] insn_o_1_925_0;
  wire  [24:0] insn_o_1_926_0;
  wire  [23:0] insn_o_1_927_0;
  wire  [23:0] insn_o_1_928_0;
  wire  [0:0] insn_o_1_929_0;
  wire  [23:0] insn_o_1_930_0;
  wire  [48:0] insn_o_1_931_0;
  wire  [0:0] insn_o_1_932_0;
  wire  [73:0] insn_o_1_933_0;
  wire  [23:0] insn_o_1_934_0;
  wire  insn_o_1_935_0;
  wire  insn_o_1_936_0;
  wire  insn_o_1_937_0;
  wire  insn_o_1_938_0;
  wire  insn_o_1_939_0;
  wire  insn_o_1_940_0;
  wire  insn_o_1_941_0;
  wire  signed [9:0] insn_o_1_942_0;
  wire  [24:0] insn_o_1_944_0;
  wire  [24:0] insn_o_1_945_0;
  wire  [23:0] insn_o_1_946_0;
  wire  [23:0] insn_o_1_947_0;
  wire  [0:0] insn_o_1_948_0;
  wire  [23:0] insn_o_1_949_0;
  wire  [48:0] insn_o_1_950_0;
  wire  [0:0] insn_o_1_951_0;
  wire  [73:0] insn_o_1_952_0;
  wire  [23:0] insn_o_1_953_0;
  wire  insn_o_1_954_0;
  wire  insn_o_1_955_0;
  wire  insn_o_1_956_0;
  wire  insn_o_1_957_0;
  wire  insn_o_1_958_0;
  wire  insn_o_1_959_0;
  wire  insn_o_1_960_0;
  wire  signed [9:0] insn_o_1_961_0;
  wire  [24:0] insn_o_1_963_0;
  wire  [24:0] insn_o_1_964_0;
  wire  [23:0] insn_o_1_965_0;
  wire  [23:0] insn_o_1_966_0;
  wire  [0:0] insn_o_1_967_0;
  wire  [23:0] insn_o_1_968_0;
  wire  [48:0] insn_o_1_969_0;
  wire  [0:0] insn_o_1_970_0;
  wire  [73:0] insn_o_1_971_0;
  wire  [23:0] insn_o_1_972_0;
  wire  insn_o_1_973_0;
  wire  insn_o_1_974_0;
  wire  insn_o_1_975_0;
  wire  insn_o_1_976_0;
  wire  insn_o_1_977_0;
  wire  insn_o_1_978_0;
  wire  insn_o_1_979_0;
  wire  signed [9:0] insn_o_1_980_0;
  wire  [24:0] insn_o_1_982_0;
  wire  [24:0] insn_o_1_983_0;
  wire  [23:0] insn_o_1_984_0;
  wire  [23:0] insn_o_1_985_0;
  wire  [0:0] insn_o_1_986_0;
  wire  [23:0] insn_o_1_987_0;
  wire  [48:0] insn_o_1_988_0;
  wire  [0:0] insn_o_1_989_0;
  wire  [73:0] insn_o_1_990_0;
  wire  [23:0] insn_o_1_991_0;
  wire  insn_o_1_992_0;
  wire  insn_o_1_993_0;
  wire  insn_o_1_994_0;
  wire  insn_o_1_995_0;
  wire  insn_o_1_996_0;
  wire  insn_o_1_997_0;
  wire  insn_o_1_998_0;
  wire  signed [9:0] insn_o_1_999_0;
  wire  [0:0] insn_o_1_1001_0;
  wire  [24:0] insn_o_1_1002_0;
  wire  [26:0] insn_o_1_1003_0;
  wire  [25:0] insn_o_1_1004_0;
  wire  [26:0] insn_o_1_1005_0;
  wire  [26:0] insn_o_1_1006_0;
  wire  [0:0] insn_o_1_1007_0;
  wire  signed [9:0] insn_o_1_1008_0;
  wire  insn_o_1_1009_0;
  wire  insn_o_1_1010_0;
  wire  insn_o_1_1011_0;
  wire  insn_o_1_1012_0;
  wire  insn_o_1_1013_0;
  wire  insn_o_1_1014_0;
  wire  insn_o_1_1015_0;
  wire  [23:0] insn_o_1_1016_0;
  wire  [0:0] insn_o_1_1017_0;
  wire  [0:0] insn_o_1_1018_0;
  wire  [0:0] insn_o_1_1019_0;
  wire  [0:0] insn_o_1_1020_0;
  wire  [0:0] insn_o_1_1021_0;
  wire  [0:0] insn_o_1_1022_0;
  wire  [0:0] insn_o_1_1023_0;
  wire  [23:0] insn_o_1_1024_0;
  wire  insn_o_1_1025_0;
  wire  [0:0] insn_o_1_1026_0;
  wire  signed [9:0] insn_o_1_1027_0;
  wire  insn_o_1_1028_0;
  wire  insn_o_1_1029_0;
  wire  insn_o_1_1030_0;
  wire  insn_o_1_1031_0;
  wire  insn_o_1_1032_0;
  wire  insn_o_1_1033_0;
  wire  insn_o_1_1034_0;
  wire  insn_o_1_1035_0;
  wire  insn_o_1_1036_0;
  wire  insn_o_1_1037_0;
  wire  [7:0] insn_o_1_1038_0;
  wire  [22:0] insn_o_1_1039_0;
  wire  [7:0] insn_o_1_1040_0;
  wire  [22:0] insn_o_1_1041_0;
  wire  [7:0] insn_o_1_1042_0;
  wire  [22:0] insn_o_1_1043_0;
  wire  insn_o_1_1044_0;
  wire  insn_o_1_1045_0;
  wire  insn_o_1_1046_0;
  wire  insn_o_1_1047_0;
  wire  insn_o_1_1048_0;
  wire  insn_o_1_1049_0;
  wire  insn_o_1_1050_0;
  wire  insn_o_1_1051_0;
  wire  insn_o_1_1052_0;
  wire  insn_o_1_1053_0;
  wire  insn_o_1_1054_0;
  wire  insn_o_1_1055_0;
  wire  insn_o_1_1056_0;
  wire  insn_o_1_1057_0;
  wire  insn_o_1_1058_0;
  wire  insn_o_1_1059_0;
  wire  insn_o_1_1060_0;
  wire  insn_o_1_1061_0;
  wire  insn_o_1_1062_0;
  wire  insn_o_1_1063_0;
  wire  insn_o_1_1064_0;
  wire  insn_o_1_1065_0;
  wire  insn_o_1_1066_0;
  wire  insn_o_1_1067_0;
  wire  insn_o_1_1068_0;
  wire  insn_o_1_1069_0;
  wire  insn_o_1_1070_0;
  wire  insn_o_1_1071_0;
  wire  insn_o_1_1072_0;
  wire  insn_o_1_1073_0;
  wire  insn_o_1_1074_0;
  wire  insn_o_1_1075_0;
  wire  insn_o_1_1076_0;
  wire  [22:0] insn_o_1_1077_0;
  wire  [7:0] insn_o_1_1078_0;
  wire  [22:0] insn_o_1_1079_0;
  wire  [7:0] insn_o_1_1080_0;
  wire  [0:0] insn_o_1_1081_0;
  wire  [22:0] insn_o_1_1082_0;
  wire  [7:0] insn_o_1_1083_0;
  wire  [31:0] insn_o_1_1084_0;
  // Insn assigns
  assign insn_o_1_4_0 = i_valid;
  assign start = insn_o_1_4_0;
  assign insn_o_1_5_0 = a_in;
  assign stage1_a_data_in = insn_o_1_5_0;
  assign insn_o_1_6_0 = stage1_a_data_in[30:23];
  assign stage1_a_exponent_in = insn_o_1_6_0;
  assign insn_o_1_7_0 = stage1_a_data_in[22:0];
  assign stage1_a_fraction_in = insn_o_1_7_0;
  assign insn_o_1_8_0 = stage1_a_data_in[31:31];
  assign stage1_a_sign_in = insn_o_1_8_0;
  assign insn_o_1_9_0 = eq_11_d0;
  assign stage1_a_exponent_zero = insn_o_1_9_0;
  assign insn_o_1_10_0 = ~stage1_a_exponent_zero;
  assign stage1_a_fraction_msb = insn_o_1_10_0;
  assign insn_o_1_11_0 = {stage1_a_fraction_msb, stage1_a_fraction_in};
  assign insn_o_1_15_0 = eq_17_d0;
  assign insn_o_1_16_0 = b_in;
  assign stage1_b_data_in = insn_o_1_16_0;
  assign insn_o_1_17_0 = stage1_b_data_in[30:23];
  assign stage1_b_exponent_in = insn_o_1_17_0;
  assign insn_o_1_18_0 = stage1_b_data_in[22:0];
  assign stage1_b_fraction_in = insn_o_1_18_0;
  assign insn_o_1_19_0 = stage1_b_data_in[31:31];
  assign stage1_b_sign_in = insn_o_1_19_0;
  assign insn_o_1_20_0 = eq_21_d0;
  assign stage1_b_exponent_zero = insn_o_1_20_0;
  assign insn_o_1_21_0 = ~stage1_b_exponent_zero;
  assign stage1_b_fraction_msb = insn_o_1_21_0;
  assign insn_o_1_22_0 = {stage1_b_fraction_msb, stage1_b_fraction_in};
  assign insn_o_1_26_0 = eq_27_d0;
  assign insn_o_1_28_0 = {2'd0, stage1_a_exponent};
  assign stage2_50_exponent_a_in = insn_o_1_28_0;
  assign insn_o_1_29_0 = sub_29_d0;
  assign stage2_50_exponent_a_d = insn_o_1_29_0;
  assign insn_o_1_30_0 = {2'd0, stage1_b_exponent};
  assign stage2_50_exponent_b_in = insn_o_1_30_0;
  assign insn_o_1_31_0 = sub_31_d0;
  assign stage2_50_exponent_b_d = insn_o_1_31_0;
  assign insn_o_1_32_0 = {25'd0, stage1_a_fraction, 25'd0};
  assign insn_o_1_34_0 = sub_34_d0;
  assign insn_o_1_35_0 = stage1_a_sign ^ stage1_b_sign;
  assign stage2_50_exponent_a_is_all_0 = stage1_a_exponent_is_all_0;
  assign insn_o_1_37_0 = eq_37_d0;
  assign stage2_50_exponent_a_is_all_1 = insn_o_1_37_0;
  assign stage2_50_fraction_a_is_all_0 = stage1_a_fraction_is_all_0;
  assign insn_o_1_39_0 = ~stage1_a_fraction_is_all_0;
  assign stage2_50_fraction_a_is_not_0 = insn_o_1_39_0;
  assign insn_o_1_40_0 = stage2_50_exponent_a_is_all_0 & stage2_50_fraction_a_is_all_0;
  assign insn_o_1_41_0 = stage2_50_exponent_a_is_all_1 & stage2_50_fraction_a_is_all_0;
  assign insn_o_1_42_0 = stage2_50_exponent_a_is_all_1 & stage2_50_fraction_a_is_not_0;
  assign stage2_50_exponent_b_is_all_0 = stage1_b_exponent_is_all_0;
  assign insn_o_1_44_0 = eq_44_d0;
  assign stage2_50_exponent_b_is_all_1 = insn_o_1_44_0;
  assign stage2_50_fraction_b_is_all_0 = stage1_b_fraction_is_all_0;
  assign insn_o_1_46_0 = ~stage1_b_fraction_is_all_0;
  assign stage2_50_fraction_b_is_not_0 = insn_o_1_46_0;
  assign insn_o_1_47_0 = stage2_50_exponent_b_is_all_0 & stage2_50_fraction_b_is_all_0;
  assign insn_o_1_48_0 = stage2_50_exponent_b_is_all_1 & stage2_50_fraction_b_is_all_0;
  assign insn_o_1_49_0 = stage2_50_exponent_b_is_all_1 & stage2_50_fraction_b_is_not_0;
  assign insn_o_1_51_0 = stage2_zi_50[73:49];
  assign stage2_49_pr = insn_o_1_51_0;
  assign insn_o_1_52_0 = sub_51_d0;
  assign stage2_49_sb = insn_o_1_52_0;
  assign insn_o_1_53_0 = stage2_49_sb[23:0];
  assign stage2_49_m0 = insn_o_1_53_0;
  assign insn_o_1_54_0 = stage2_49_pr[23:0];
  assign stage2_49_m1 = insn_o_1_54_0;
  assign insn_o_1_55_0 = stage2_49_sb[24:24];
  assign stage2_49_ms = insn_o_1_55_0;
  assign insn_o_1_56_0 = stage2_49_ms ? stage2_49_m1 : stage2_49_m0;
  assign stage2_49_mx = insn_o_1_56_0;
  assign insn_o_1_57_0 = stage2_zi_50[48:0];
  assign stage2_49_zl = insn_o_1_57_0;
  assign insn_o_1_58_0 = ~stage2_49_ms;
  assign stage2_49_zb = insn_o_1_58_0;
  assign insn_o_1_59_0 = {stage2_49_mx, stage2_49_zl, stage2_49_zb};
  assign insn_o_1_70_0 = stage2_zi_49[73:49];
  assign stage2_48_pr = insn_o_1_70_0;
  assign insn_o_1_71_0 = sub_69_d0;
  assign stage2_48_sb = insn_o_1_71_0;
  assign insn_o_1_72_0 = stage2_48_sb[23:0];
  assign stage2_48_m0 = insn_o_1_72_0;
  assign insn_o_1_73_0 = stage2_48_pr[23:0];
  assign stage2_48_m1 = insn_o_1_73_0;
  assign insn_o_1_74_0 = stage2_48_sb[24:24];
  assign stage2_48_ms = insn_o_1_74_0;
  assign insn_o_1_75_0 = stage2_48_ms ? stage2_48_m1 : stage2_48_m0;
  assign stage2_48_mx = insn_o_1_75_0;
  assign insn_o_1_76_0 = stage2_zi_49[48:0];
  assign stage2_48_zl = insn_o_1_76_0;
  assign insn_o_1_77_0 = ~stage2_48_ms;
  assign stage2_48_zb = insn_o_1_77_0;
  assign insn_o_1_78_0 = {stage2_48_mx, stage2_48_zl, stage2_48_zb};
  assign insn_o_1_89_0 = stage2_zi_48[73:49];
  assign stage2_47_pr = insn_o_1_89_0;
  assign insn_o_1_90_0 = sub_87_d0;
  assign stage2_47_sb = insn_o_1_90_0;
  assign insn_o_1_91_0 = stage2_47_sb[23:0];
  assign stage2_47_m0 = insn_o_1_91_0;
  assign insn_o_1_92_0 = stage2_47_pr[23:0];
  assign stage2_47_m1 = insn_o_1_92_0;
  assign insn_o_1_93_0 = stage2_47_sb[24:24];
  assign stage2_47_ms = insn_o_1_93_0;
  assign insn_o_1_94_0 = stage2_47_ms ? stage2_47_m1 : stage2_47_m0;
  assign stage2_47_mx = insn_o_1_94_0;
  assign insn_o_1_95_0 = stage2_zi_48[48:0];
  assign stage2_47_zl = insn_o_1_95_0;
  assign insn_o_1_96_0 = ~stage2_47_ms;
  assign stage2_47_zb = insn_o_1_96_0;
  assign insn_o_1_97_0 = {stage2_47_mx, stage2_47_zl, stage2_47_zb};
  assign insn_o_1_108_0 = stage2_zi_47[73:49];
  assign stage2_46_pr = insn_o_1_108_0;
  assign insn_o_1_109_0 = sub_105_d0;
  assign stage2_46_sb = insn_o_1_109_0;
  assign insn_o_1_110_0 = stage2_46_sb[23:0];
  assign stage2_46_m0 = insn_o_1_110_0;
  assign insn_o_1_111_0 = stage2_46_pr[23:0];
  assign stage2_46_m1 = insn_o_1_111_0;
  assign insn_o_1_112_0 = stage2_46_sb[24:24];
  assign stage2_46_ms = insn_o_1_112_0;
  assign insn_o_1_113_0 = stage2_46_ms ? stage2_46_m1 : stage2_46_m0;
  assign stage2_46_mx = insn_o_1_113_0;
  assign insn_o_1_114_0 = stage2_zi_47[48:0];
  assign stage2_46_zl = insn_o_1_114_0;
  assign insn_o_1_115_0 = ~stage2_46_ms;
  assign stage2_46_zb = insn_o_1_115_0;
  assign insn_o_1_116_0 = {stage2_46_mx, stage2_46_zl, stage2_46_zb};
  assign insn_o_1_127_0 = stage2_zi_46[73:49];
  assign stage2_45_pr = insn_o_1_127_0;
  assign insn_o_1_128_0 = sub_123_d0;
  assign stage2_45_sb = insn_o_1_128_0;
  assign insn_o_1_129_0 = stage2_45_sb[23:0];
  assign stage2_45_m0 = insn_o_1_129_0;
  assign insn_o_1_130_0 = stage2_45_pr[23:0];
  assign stage2_45_m1 = insn_o_1_130_0;
  assign insn_o_1_131_0 = stage2_45_sb[24:24];
  assign stage2_45_ms = insn_o_1_131_0;
  assign insn_o_1_132_0 = stage2_45_ms ? stage2_45_m1 : stage2_45_m0;
  assign stage2_45_mx = insn_o_1_132_0;
  assign insn_o_1_133_0 = stage2_zi_46[48:0];
  assign stage2_45_zl = insn_o_1_133_0;
  assign insn_o_1_134_0 = ~stage2_45_ms;
  assign stage2_45_zb = insn_o_1_134_0;
  assign insn_o_1_135_0 = {stage2_45_mx, stage2_45_zl, stage2_45_zb};
  assign insn_o_1_146_0 = stage2_zi_45[73:49];
  assign stage2_44_pr = insn_o_1_146_0;
  assign insn_o_1_147_0 = sub_141_d0;
  assign stage2_44_sb = insn_o_1_147_0;
  assign insn_o_1_148_0 = stage2_44_sb[23:0];
  assign stage2_44_m0 = insn_o_1_148_0;
  assign insn_o_1_149_0 = stage2_44_pr[23:0];
  assign stage2_44_m1 = insn_o_1_149_0;
  assign insn_o_1_150_0 = stage2_44_sb[24:24];
  assign stage2_44_ms = insn_o_1_150_0;
  assign insn_o_1_151_0 = stage2_44_ms ? stage2_44_m1 : stage2_44_m0;
  assign stage2_44_mx = insn_o_1_151_0;
  assign insn_o_1_152_0 = stage2_zi_45[48:0];
  assign stage2_44_zl = insn_o_1_152_0;
  assign insn_o_1_153_0 = ~stage2_44_ms;
  assign stage2_44_zb = insn_o_1_153_0;
  assign insn_o_1_154_0 = {stage2_44_mx, stage2_44_zl, stage2_44_zb};
  assign insn_o_1_165_0 = stage2_zi_44[73:49];
  assign stage2_43_pr = insn_o_1_165_0;
  assign insn_o_1_166_0 = sub_159_d0;
  assign stage2_43_sb = insn_o_1_166_0;
  assign insn_o_1_167_0 = stage2_43_sb[23:0];
  assign stage2_43_m0 = insn_o_1_167_0;
  assign insn_o_1_168_0 = stage2_43_pr[23:0];
  assign stage2_43_m1 = insn_o_1_168_0;
  assign insn_o_1_169_0 = stage2_43_sb[24:24];
  assign stage2_43_ms = insn_o_1_169_0;
  assign insn_o_1_170_0 = stage2_43_ms ? stage2_43_m1 : stage2_43_m0;
  assign stage2_43_mx = insn_o_1_170_0;
  assign insn_o_1_171_0 = stage2_zi_44[48:0];
  assign stage2_43_zl = insn_o_1_171_0;
  assign insn_o_1_172_0 = ~stage2_43_ms;
  assign stage2_43_zb = insn_o_1_172_0;
  assign insn_o_1_173_0 = {stage2_43_mx, stage2_43_zl, stage2_43_zb};
  assign insn_o_1_184_0 = stage2_zi_43[73:49];
  assign stage2_42_pr = insn_o_1_184_0;
  assign insn_o_1_185_0 = sub_177_d0;
  assign stage2_42_sb = insn_o_1_185_0;
  assign insn_o_1_186_0 = stage2_42_sb[23:0];
  assign stage2_42_m0 = insn_o_1_186_0;
  assign insn_o_1_187_0 = stage2_42_pr[23:0];
  assign stage2_42_m1 = insn_o_1_187_0;
  assign insn_o_1_188_0 = stage2_42_sb[24:24];
  assign stage2_42_ms = insn_o_1_188_0;
  assign insn_o_1_189_0 = stage2_42_ms ? stage2_42_m1 : stage2_42_m0;
  assign stage2_42_mx = insn_o_1_189_0;
  assign insn_o_1_190_0 = stage2_zi_43[48:0];
  assign stage2_42_zl = insn_o_1_190_0;
  assign insn_o_1_191_0 = ~stage2_42_ms;
  assign stage2_42_zb = insn_o_1_191_0;
  assign insn_o_1_192_0 = {stage2_42_mx, stage2_42_zl, stage2_42_zb};
  assign insn_o_1_203_0 = stage2_zi_42[73:49];
  assign stage2_41_pr = insn_o_1_203_0;
  assign insn_o_1_204_0 = sub_195_d0;
  assign stage2_41_sb = insn_o_1_204_0;
  assign insn_o_1_205_0 = stage2_41_sb[23:0];
  assign stage2_41_m0 = insn_o_1_205_0;
  assign insn_o_1_206_0 = stage2_41_pr[23:0];
  assign stage2_41_m1 = insn_o_1_206_0;
  assign insn_o_1_207_0 = stage2_41_sb[24:24];
  assign stage2_41_ms = insn_o_1_207_0;
  assign insn_o_1_208_0 = stage2_41_ms ? stage2_41_m1 : stage2_41_m0;
  assign stage2_41_mx = insn_o_1_208_0;
  assign insn_o_1_209_0 = stage2_zi_42[48:0];
  assign stage2_41_zl = insn_o_1_209_0;
  assign insn_o_1_210_0 = ~stage2_41_ms;
  assign stage2_41_zb = insn_o_1_210_0;
  assign insn_o_1_211_0 = {stage2_41_mx, stage2_41_zl, stage2_41_zb};
  assign insn_o_1_222_0 = stage2_zi_41[73:49];
  assign stage2_40_pr = insn_o_1_222_0;
  assign insn_o_1_223_0 = sub_213_d0;
  assign stage2_40_sb = insn_o_1_223_0;
  assign insn_o_1_224_0 = stage2_40_sb[23:0];
  assign stage2_40_m0 = insn_o_1_224_0;
  assign insn_o_1_225_0 = stage2_40_pr[23:0];
  assign stage2_40_m1 = insn_o_1_225_0;
  assign insn_o_1_226_0 = stage2_40_sb[24:24];
  assign stage2_40_ms = insn_o_1_226_0;
  assign insn_o_1_227_0 = stage2_40_ms ? stage2_40_m1 : stage2_40_m0;
  assign stage2_40_mx = insn_o_1_227_0;
  assign insn_o_1_228_0 = stage2_zi_41[48:0];
  assign stage2_40_zl = insn_o_1_228_0;
  assign insn_o_1_229_0 = ~stage2_40_ms;
  assign stage2_40_zb = insn_o_1_229_0;
  assign insn_o_1_230_0 = {stage2_40_mx, stage2_40_zl, stage2_40_zb};
  assign insn_o_1_241_0 = stage2_zi_40[73:49];
  assign stage2_39_pr = insn_o_1_241_0;
  assign insn_o_1_242_0 = sub_231_d0;
  assign stage2_39_sb = insn_o_1_242_0;
  assign insn_o_1_243_0 = stage2_39_sb[23:0];
  assign stage2_39_m0 = insn_o_1_243_0;
  assign insn_o_1_244_0 = stage2_39_pr[23:0];
  assign stage2_39_m1 = insn_o_1_244_0;
  assign insn_o_1_245_0 = stage2_39_sb[24:24];
  assign stage2_39_ms = insn_o_1_245_0;
  assign insn_o_1_246_0 = stage2_39_ms ? stage2_39_m1 : stage2_39_m0;
  assign stage2_39_mx = insn_o_1_246_0;
  assign insn_o_1_247_0 = stage2_zi_40[48:0];
  assign stage2_39_zl = insn_o_1_247_0;
  assign insn_o_1_248_0 = ~stage2_39_ms;
  assign stage2_39_zb = insn_o_1_248_0;
  assign insn_o_1_249_0 = {stage2_39_mx, stage2_39_zl, stage2_39_zb};
  assign insn_o_1_260_0 = stage2_zi_39[73:49];
  assign stage2_38_pr = insn_o_1_260_0;
  assign insn_o_1_261_0 = sub_249_d0;
  assign stage2_38_sb = insn_o_1_261_0;
  assign insn_o_1_262_0 = stage2_38_sb[23:0];
  assign stage2_38_m0 = insn_o_1_262_0;
  assign insn_o_1_263_0 = stage2_38_pr[23:0];
  assign stage2_38_m1 = insn_o_1_263_0;
  assign insn_o_1_264_0 = stage2_38_sb[24:24];
  assign stage2_38_ms = insn_o_1_264_0;
  assign insn_o_1_265_0 = stage2_38_ms ? stage2_38_m1 : stage2_38_m0;
  assign stage2_38_mx = insn_o_1_265_0;
  assign insn_o_1_266_0 = stage2_zi_39[48:0];
  assign stage2_38_zl = insn_o_1_266_0;
  assign insn_o_1_267_0 = ~stage2_38_ms;
  assign stage2_38_zb = insn_o_1_267_0;
  assign insn_o_1_268_0 = {stage2_38_mx, stage2_38_zl, stage2_38_zb};
  assign insn_o_1_279_0 = stage2_zi_38[73:49];
  assign stage2_37_pr = insn_o_1_279_0;
  assign insn_o_1_280_0 = sub_267_d0;
  assign stage2_37_sb = insn_o_1_280_0;
  assign insn_o_1_281_0 = stage2_37_sb[23:0];
  assign stage2_37_m0 = insn_o_1_281_0;
  assign insn_o_1_282_0 = stage2_37_pr[23:0];
  assign stage2_37_m1 = insn_o_1_282_0;
  assign insn_o_1_283_0 = stage2_37_sb[24:24];
  assign stage2_37_ms = insn_o_1_283_0;
  assign insn_o_1_284_0 = stage2_37_ms ? stage2_37_m1 : stage2_37_m0;
  assign stage2_37_mx = insn_o_1_284_0;
  assign insn_o_1_285_0 = stage2_zi_38[48:0];
  assign stage2_37_zl = insn_o_1_285_0;
  assign insn_o_1_286_0 = ~stage2_37_ms;
  assign stage2_37_zb = insn_o_1_286_0;
  assign insn_o_1_287_0 = {stage2_37_mx, stage2_37_zl, stage2_37_zb};
  assign insn_o_1_298_0 = stage2_zi_37[73:49];
  assign stage2_36_pr = insn_o_1_298_0;
  assign insn_o_1_299_0 = sub_285_d0;
  assign stage2_36_sb = insn_o_1_299_0;
  assign insn_o_1_300_0 = stage2_36_sb[23:0];
  assign stage2_36_m0 = insn_o_1_300_0;
  assign insn_o_1_301_0 = stage2_36_pr[23:0];
  assign stage2_36_m1 = insn_o_1_301_0;
  assign insn_o_1_302_0 = stage2_36_sb[24:24];
  assign stage2_36_ms = insn_o_1_302_0;
  assign insn_o_1_303_0 = stage2_36_ms ? stage2_36_m1 : stage2_36_m0;
  assign stage2_36_mx = insn_o_1_303_0;
  assign insn_o_1_304_0 = stage2_zi_37[48:0];
  assign stage2_36_zl = insn_o_1_304_0;
  assign insn_o_1_305_0 = ~stage2_36_ms;
  assign stage2_36_zb = insn_o_1_305_0;
  assign insn_o_1_306_0 = {stage2_36_mx, stage2_36_zl, stage2_36_zb};
  assign insn_o_1_317_0 = stage2_zi_36[73:49];
  assign stage2_35_pr = insn_o_1_317_0;
  assign insn_o_1_318_0 = sub_303_d0;
  assign stage2_35_sb = insn_o_1_318_0;
  assign insn_o_1_319_0 = stage2_35_sb[23:0];
  assign stage2_35_m0 = insn_o_1_319_0;
  assign insn_o_1_320_0 = stage2_35_pr[23:0];
  assign stage2_35_m1 = insn_o_1_320_0;
  assign insn_o_1_321_0 = stage2_35_sb[24:24];
  assign stage2_35_ms = insn_o_1_321_0;
  assign insn_o_1_322_0 = stage2_35_ms ? stage2_35_m1 : stage2_35_m0;
  assign stage2_35_mx = insn_o_1_322_0;
  assign insn_o_1_323_0 = stage2_zi_36[48:0];
  assign stage2_35_zl = insn_o_1_323_0;
  assign insn_o_1_324_0 = ~stage2_35_ms;
  assign stage2_35_zb = insn_o_1_324_0;
  assign insn_o_1_325_0 = {stage2_35_mx, stage2_35_zl, stage2_35_zb};
  assign insn_o_1_336_0 = stage2_zi_35[73:49];
  assign stage2_34_pr = insn_o_1_336_0;
  assign insn_o_1_337_0 = sub_321_d0;
  assign stage2_34_sb = insn_o_1_337_0;
  assign insn_o_1_338_0 = stage2_34_sb[23:0];
  assign stage2_34_m0 = insn_o_1_338_0;
  assign insn_o_1_339_0 = stage2_34_pr[23:0];
  assign stage2_34_m1 = insn_o_1_339_0;
  assign insn_o_1_340_0 = stage2_34_sb[24:24];
  assign stage2_34_ms = insn_o_1_340_0;
  assign insn_o_1_341_0 = stage2_34_ms ? stage2_34_m1 : stage2_34_m0;
  assign stage2_34_mx = insn_o_1_341_0;
  assign insn_o_1_342_0 = stage2_zi_35[48:0];
  assign stage2_34_zl = insn_o_1_342_0;
  assign insn_o_1_343_0 = ~stage2_34_ms;
  assign stage2_34_zb = insn_o_1_343_0;
  assign insn_o_1_344_0 = {stage2_34_mx, stage2_34_zl, stage2_34_zb};
  assign insn_o_1_355_0 = stage2_zi_34[73:49];
  assign stage2_33_pr = insn_o_1_355_0;
  assign insn_o_1_356_0 = sub_339_d0;
  assign stage2_33_sb = insn_o_1_356_0;
  assign insn_o_1_357_0 = stage2_33_sb[23:0];
  assign stage2_33_m0 = insn_o_1_357_0;
  assign insn_o_1_358_0 = stage2_33_pr[23:0];
  assign stage2_33_m1 = insn_o_1_358_0;
  assign insn_o_1_359_0 = stage2_33_sb[24:24];
  assign stage2_33_ms = insn_o_1_359_0;
  assign insn_o_1_360_0 = stage2_33_ms ? stage2_33_m1 : stage2_33_m0;
  assign stage2_33_mx = insn_o_1_360_0;
  assign insn_o_1_361_0 = stage2_zi_34[48:0];
  assign stage2_33_zl = insn_o_1_361_0;
  assign insn_o_1_362_0 = ~stage2_33_ms;
  assign stage2_33_zb = insn_o_1_362_0;
  assign insn_o_1_363_0 = {stage2_33_mx, stage2_33_zl, stage2_33_zb};
  assign insn_o_1_374_0 = stage2_zi_33[73:49];
  assign stage2_32_pr = insn_o_1_374_0;
  assign insn_o_1_375_0 = sub_357_d0;
  assign stage2_32_sb = insn_o_1_375_0;
  assign insn_o_1_376_0 = stage2_32_sb[23:0];
  assign stage2_32_m0 = insn_o_1_376_0;
  assign insn_o_1_377_0 = stage2_32_pr[23:0];
  assign stage2_32_m1 = insn_o_1_377_0;
  assign insn_o_1_378_0 = stage2_32_sb[24:24];
  assign stage2_32_ms = insn_o_1_378_0;
  assign insn_o_1_379_0 = stage2_32_ms ? stage2_32_m1 : stage2_32_m0;
  assign stage2_32_mx = insn_o_1_379_0;
  assign insn_o_1_380_0 = stage2_zi_33[48:0];
  assign stage2_32_zl = insn_o_1_380_0;
  assign insn_o_1_381_0 = ~stage2_32_ms;
  assign stage2_32_zb = insn_o_1_381_0;
  assign insn_o_1_382_0 = {stage2_32_mx, stage2_32_zl, stage2_32_zb};
  assign insn_o_1_393_0 = stage2_zi_32[73:49];
  assign stage2_31_pr = insn_o_1_393_0;
  assign insn_o_1_394_0 = sub_375_d0;
  assign stage2_31_sb = insn_o_1_394_0;
  assign insn_o_1_395_0 = stage2_31_sb[23:0];
  assign stage2_31_m0 = insn_o_1_395_0;
  assign insn_o_1_396_0 = stage2_31_pr[23:0];
  assign stage2_31_m1 = insn_o_1_396_0;
  assign insn_o_1_397_0 = stage2_31_sb[24:24];
  assign stage2_31_ms = insn_o_1_397_0;
  assign insn_o_1_398_0 = stage2_31_ms ? stage2_31_m1 : stage2_31_m0;
  assign stage2_31_mx = insn_o_1_398_0;
  assign insn_o_1_399_0 = stage2_zi_32[48:0];
  assign stage2_31_zl = insn_o_1_399_0;
  assign insn_o_1_400_0 = ~stage2_31_ms;
  assign stage2_31_zb = insn_o_1_400_0;
  assign insn_o_1_401_0 = {stage2_31_mx, stage2_31_zl, stage2_31_zb};
  assign insn_o_1_412_0 = stage2_zi_31[73:49];
  assign stage2_30_pr = insn_o_1_412_0;
  assign insn_o_1_413_0 = sub_393_d0;
  assign stage2_30_sb = insn_o_1_413_0;
  assign insn_o_1_414_0 = stage2_30_sb[23:0];
  assign stage2_30_m0 = insn_o_1_414_0;
  assign insn_o_1_415_0 = stage2_30_pr[23:0];
  assign stage2_30_m1 = insn_o_1_415_0;
  assign insn_o_1_416_0 = stage2_30_sb[24:24];
  assign stage2_30_ms = insn_o_1_416_0;
  assign insn_o_1_417_0 = stage2_30_ms ? stage2_30_m1 : stage2_30_m0;
  assign stage2_30_mx = insn_o_1_417_0;
  assign insn_o_1_418_0 = stage2_zi_31[48:0];
  assign stage2_30_zl = insn_o_1_418_0;
  assign insn_o_1_419_0 = ~stage2_30_ms;
  assign stage2_30_zb = insn_o_1_419_0;
  assign insn_o_1_420_0 = {stage2_30_mx, stage2_30_zl, stage2_30_zb};
  assign insn_o_1_431_0 = stage2_zi_30[73:49];
  assign stage2_29_pr = insn_o_1_431_0;
  assign insn_o_1_432_0 = sub_411_d0;
  assign stage2_29_sb = insn_o_1_432_0;
  assign insn_o_1_433_0 = stage2_29_sb[23:0];
  assign stage2_29_m0 = insn_o_1_433_0;
  assign insn_o_1_434_0 = stage2_29_pr[23:0];
  assign stage2_29_m1 = insn_o_1_434_0;
  assign insn_o_1_435_0 = stage2_29_sb[24:24];
  assign stage2_29_ms = insn_o_1_435_0;
  assign insn_o_1_436_0 = stage2_29_ms ? stage2_29_m1 : stage2_29_m0;
  assign stage2_29_mx = insn_o_1_436_0;
  assign insn_o_1_437_0 = stage2_zi_30[48:0];
  assign stage2_29_zl = insn_o_1_437_0;
  assign insn_o_1_438_0 = ~stage2_29_ms;
  assign stage2_29_zb = insn_o_1_438_0;
  assign insn_o_1_439_0 = {stage2_29_mx, stage2_29_zl, stage2_29_zb};
  assign insn_o_1_450_0 = stage2_zi_29[73:49];
  assign stage2_28_pr = insn_o_1_450_0;
  assign insn_o_1_451_0 = sub_429_d0;
  assign stage2_28_sb = insn_o_1_451_0;
  assign insn_o_1_452_0 = stage2_28_sb[23:0];
  assign stage2_28_m0 = insn_o_1_452_0;
  assign insn_o_1_453_0 = stage2_28_pr[23:0];
  assign stage2_28_m1 = insn_o_1_453_0;
  assign insn_o_1_454_0 = stage2_28_sb[24:24];
  assign stage2_28_ms = insn_o_1_454_0;
  assign insn_o_1_455_0 = stage2_28_ms ? stage2_28_m1 : stage2_28_m0;
  assign stage2_28_mx = insn_o_1_455_0;
  assign insn_o_1_456_0 = stage2_zi_29[48:0];
  assign stage2_28_zl = insn_o_1_456_0;
  assign insn_o_1_457_0 = ~stage2_28_ms;
  assign stage2_28_zb = insn_o_1_457_0;
  assign insn_o_1_458_0 = {stage2_28_mx, stage2_28_zl, stage2_28_zb};
  assign insn_o_1_469_0 = stage2_zi_28[73:49];
  assign stage2_27_pr = insn_o_1_469_0;
  assign insn_o_1_470_0 = sub_447_d0;
  assign stage2_27_sb = insn_o_1_470_0;
  assign insn_o_1_471_0 = stage2_27_sb[23:0];
  assign stage2_27_m0 = insn_o_1_471_0;
  assign insn_o_1_472_0 = stage2_27_pr[23:0];
  assign stage2_27_m1 = insn_o_1_472_0;
  assign insn_o_1_473_0 = stage2_27_sb[24:24];
  assign stage2_27_ms = insn_o_1_473_0;
  assign insn_o_1_474_0 = stage2_27_ms ? stage2_27_m1 : stage2_27_m0;
  assign stage2_27_mx = insn_o_1_474_0;
  assign insn_o_1_475_0 = stage2_zi_28[48:0];
  assign stage2_27_zl = insn_o_1_475_0;
  assign insn_o_1_476_0 = ~stage2_27_ms;
  assign stage2_27_zb = insn_o_1_476_0;
  assign insn_o_1_477_0 = {stage2_27_mx, stage2_27_zl, stage2_27_zb};
  assign insn_o_1_488_0 = stage2_zi_27[73:49];
  assign stage2_26_pr = insn_o_1_488_0;
  assign insn_o_1_489_0 = sub_465_d0;
  assign stage2_26_sb = insn_o_1_489_0;
  assign insn_o_1_490_0 = stage2_26_sb[23:0];
  assign stage2_26_m0 = insn_o_1_490_0;
  assign insn_o_1_491_0 = stage2_26_pr[23:0];
  assign stage2_26_m1 = insn_o_1_491_0;
  assign insn_o_1_492_0 = stage2_26_sb[24:24];
  assign stage2_26_ms = insn_o_1_492_0;
  assign insn_o_1_493_0 = stage2_26_ms ? stage2_26_m1 : stage2_26_m0;
  assign stage2_26_mx = insn_o_1_493_0;
  assign insn_o_1_494_0 = stage2_zi_27[48:0];
  assign stage2_26_zl = insn_o_1_494_0;
  assign insn_o_1_495_0 = ~stage2_26_ms;
  assign stage2_26_zb = insn_o_1_495_0;
  assign insn_o_1_496_0 = {stage2_26_mx, stage2_26_zl, stage2_26_zb};
  assign insn_o_1_507_0 = stage2_zi_26[73:49];
  assign stage2_25_pr = insn_o_1_507_0;
  assign insn_o_1_508_0 = sub_483_d0;
  assign stage2_25_sb = insn_o_1_508_0;
  assign insn_o_1_509_0 = stage2_25_sb[23:0];
  assign stage2_25_m0 = insn_o_1_509_0;
  assign insn_o_1_510_0 = stage2_25_pr[23:0];
  assign stage2_25_m1 = insn_o_1_510_0;
  assign insn_o_1_511_0 = stage2_25_sb[24:24];
  assign stage2_25_ms = insn_o_1_511_0;
  assign insn_o_1_512_0 = stage2_25_ms ? stage2_25_m1 : stage2_25_m0;
  assign stage2_25_mx = insn_o_1_512_0;
  assign insn_o_1_513_0 = stage2_zi_26[48:0];
  assign stage2_25_zl = insn_o_1_513_0;
  assign insn_o_1_514_0 = ~stage2_25_ms;
  assign stage2_25_zb = insn_o_1_514_0;
  assign insn_o_1_515_0 = {stage2_25_mx, stage2_25_zl, stage2_25_zb};
  assign insn_o_1_526_0 = stage2_zi_25[73:49];
  assign stage2_24_pr = insn_o_1_526_0;
  assign insn_o_1_527_0 = sub_501_d0;
  assign stage2_24_sb = insn_o_1_527_0;
  assign insn_o_1_528_0 = stage2_24_sb[23:0];
  assign stage2_24_m0 = insn_o_1_528_0;
  assign insn_o_1_529_0 = stage2_24_pr[23:0];
  assign stage2_24_m1 = insn_o_1_529_0;
  assign insn_o_1_530_0 = stage2_24_sb[24:24];
  assign stage2_24_ms = insn_o_1_530_0;
  assign insn_o_1_531_0 = stage2_24_ms ? stage2_24_m1 : stage2_24_m0;
  assign stage2_24_mx = insn_o_1_531_0;
  assign insn_o_1_532_0 = stage2_zi_25[48:0];
  assign stage2_24_zl = insn_o_1_532_0;
  assign insn_o_1_533_0 = ~stage2_24_ms;
  assign stage2_24_zb = insn_o_1_533_0;
  assign insn_o_1_534_0 = {stage2_24_mx, stage2_24_zl, stage2_24_zb};
  assign insn_o_1_545_0 = stage2_zi_24[73:49];
  assign stage2_23_pr = insn_o_1_545_0;
  assign insn_o_1_546_0 = sub_519_d0;
  assign stage2_23_sb = insn_o_1_546_0;
  assign insn_o_1_547_0 = stage2_23_sb[23:0];
  assign stage2_23_m0 = insn_o_1_547_0;
  assign insn_o_1_548_0 = stage2_23_pr[23:0];
  assign stage2_23_m1 = insn_o_1_548_0;
  assign insn_o_1_549_0 = stage2_23_sb[24:24];
  assign stage2_23_ms = insn_o_1_549_0;
  assign insn_o_1_550_0 = stage2_23_ms ? stage2_23_m1 : stage2_23_m0;
  assign stage2_23_mx = insn_o_1_550_0;
  assign insn_o_1_551_0 = stage2_zi_24[48:0];
  assign stage2_23_zl = insn_o_1_551_0;
  assign insn_o_1_552_0 = ~stage2_23_ms;
  assign stage2_23_zb = insn_o_1_552_0;
  assign insn_o_1_553_0 = {stage2_23_mx, stage2_23_zl, stage2_23_zb};
  assign insn_o_1_564_0 = stage2_zi_23[73:49];
  assign stage2_22_pr = insn_o_1_564_0;
  assign insn_o_1_565_0 = sub_537_d0;
  assign stage2_22_sb = insn_o_1_565_0;
  assign insn_o_1_566_0 = stage2_22_sb[23:0];
  assign stage2_22_m0 = insn_o_1_566_0;
  assign insn_o_1_567_0 = stage2_22_pr[23:0];
  assign stage2_22_m1 = insn_o_1_567_0;
  assign insn_o_1_568_0 = stage2_22_sb[24:24];
  assign stage2_22_ms = insn_o_1_568_0;
  assign insn_o_1_569_0 = stage2_22_ms ? stage2_22_m1 : stage2_22_m0;
  assign stage2_22_mx = insn_o_1_569_0;
  assign insn_o_1_570_0 = stage2_zi_23[48:0];
  assign stage2_22_zl = insn_o_1_570_0;
  assign insn_o_1_571_0 = ~stage2_22_ms;
  assign stage2_22_zb = insn_o_1_571_0;
  assign insn_o_1_572_0 = {stage2_22_mx, stage2_22_zl, stage2_22_zb};
  assign insn_o_1_583_0 = stage2_zi_22[73:49];
  assign stage2_21_pr = insn_o_1_583_0;
  assign insn_o_1_584_0 = sub_555_d0;
  assign stage2_21_sb = insn_o_1_584_0;
  assign insn_o_1_585_0 = stage2_21_sb[23:0];
  assign stage2_21_m0 = insn_o_1_585_0;
  assign insn_o_1_586_0 = stage2_21_pr[23:0];
  assign stage2_21_m1 = insn_o_1_586_0;
  assign insn_o_1_587_0 = stage2_21_sb[24:24];
  assign stage2_21_ms = insn_o_1_587_0;
  assign insn_o_1_588_0 = stage2_21_ms ? stage2_21_m1 : stage2_21_m0;
  assign stage2_21_mx = insn_o_1_588_0;
  assign insn_o_1_589_0 = stage2_zi_22[48:0];
  assign stage2_21_zl = insn_o_1_589_0;
  assign insn_o_1_590_0 = ~stage2_21_ms;
  assign stage2_21_zb = insn_o_1_590_0;
  assign insn_o_1_591_0 = {stage2_21_mx, stage2_21_zl, stage2_21_zb};
  assign insn_o_1_602_0 = stage2_zi_21[73:49];
  assign stage2_20_pr = insn_o_1_602_0;
  assign insn_o_1_603_0 = sub_573_d0;
  assign stage2_20_sb = insn_o_1_603_0;
  assign insn_o_1_604_0 = stage2_20_sb[23:0];
  assign stage2_20_m0 = insn_o_1_604_0;
  assign insn_o_1_605_0 = stage2_20_pr[23:0];
  assign stage2_20_m1 = insn_o_1_605_0;
  assign insn_o_1_606_0 = stage2_20_sb[24:24];
  assign stage2_20_ms = insn_o_1_606_0;
  assign insn_o_1_607_0 = stage2_20_ms ? stage2_20_m1 : stage2_20_m0;
  assign stage2_20_mx = insn_o_1_607_0;
  assign insn_o_1_608_0 = stage2_zi_21[48:0];
  assign stage2_20_zl = insn_o_1_608_0;
  assign insn_o_1_609_0 = ~stage2_20_ms;
  assign stage2_20_zb = insn_o_1_609_0;
  assign insn_o_1_610_0 = {stage2_20_mx, stage2_20_zl, stage2_20_zb};
  assign insn_o_1_621_0 = stage2_zi_20[73:49];
  assign stage2_19_pr = insn_o_1_621_0;
  assign insn_o_1_622_0 = sub_591_d0;
  assign stage2_19_sb = insn_o_1_622_0;
  assign insn_o_1_623_0 = stage2_19_sb[23:0];
  assign stage2_19_m0 = insn_o_1_623_0;
  assign insn_o_1_624_0 = stage2_19_pr[23:0];
  assign stage2_19_m1 = insn_o_1_624_0;
  assign insn_o_1_625_0 = stage2_19_sb[24:24];
  assign stage2_19_ms = insn_o_1_625_0;
  assign insn_o_1_626_0 = stage2_19_ms ? stage2_19_m1 : stage2_19_m0;
  assign stage2_19_mx = insn_o_1_626_0;
  assign insn_o_1_627_0 = stage2_zi_20[48:0];
  assign stage2_19_zl = insn_o_1_627_0;
  assign insn_o_1_628_0 = ~stage2_19_ms;
  assign stage2_19_zb = insn_o_1_628_0;
  assign insn_o_1_629_0 = {stage2_19_mx, stage2_19_zl, stage2_19_zb};
  assign insn_o_1_640_0 = stage2_zi_19[73:49];
  assign stage2_18_pr = insn_o_1_640_0;
  assign insn_o_1_641_0 = sub_609_d0;
  assign stage2_18_sb = insn_o_1_641_0;
  assign insn_o_1_642_0 = stage2_18_sb[23:0];
  assign stage2_18_m0 = insn_o_1_642_0;
  assign insn_o_1_643_0 = stage2_18_pr[23:0];
  assign stage2_18_m1 = insn_o_1_643_0;
  assign insn_o_1_644_0 = stage2_18_sb[24:24];
  assign stage2_18_ms = insn_o_1_644_0;
  assign insn_o_1_645_0 = stage2_18_ms ? stage2_18_m1 : stage2_18_m0;
  assign stage2_18_mx = insn_o_1_645_0;
  assign insn_o_1_646_0 = stage2_zi_19[48:0];
  assign stage2_18_zl = insn_o_1_646_0;
  assign insn_o_1_647_0 = ~stage2_18_ms;
  assign stage2_18_zb = insn_o_1_647_0;
  assign insn_o_1_648_0 = {stage2_18_mx, stage2_18_zl, stage2_18_zb};
  assign insn_o_1_659_0 = stage2_zi_18[73:49];
  assign stage2_17_pr = insn_o_1_659_0;
  assign insn_o_1_660_0 = sub_627_d0;
  assign stage2_17_sb = insn_o_1_660_0;
  assign insn_o_1_661_0 = stage2_17_sb[23:0];
  assign stage2_17_m0 = insn_o_1_661_0;
  assign insn_o_1_662_0 = stage2_17_pr[23:0];
  assign stage2_17_m1 = insn_o_1_662_0;
  assign insn_o_1_663_0 = stage2_17_sb[24:24];
  assign stage2_17_ms = insn_o_1_663_0;
  assign insn_o_1_664_0 = stage2_17_ms ? stage2_17_m1 : stage2_17_m0;
  assign stage2_17_mx = insn_o_1_664_0;
  assign insn_o_1_665_0 = stage2_zi_18[48:0];
  assign stage2_17_zl = insn_o_1_665_0;
  assign insn_o_1_666_0 = ~stage2_17_ms;
  assign stage2_17_zb = insn_o_1_666_0;
  assign insn_o_1_667_0 = {stage2_17_mx, stage2_17_zl, stage2_17_zb};
  assign insn_o_1_678_0 = stage2_zi_17[73:49];
  assign stage2_16_pr = insn_o_1_678_0;
  assign insn_o_1_679_0 = sub_645_d0;
  assign stage2_16_sb = insn_o_1_679_0;
  assign insn_o_1_680_0 = stage2_16_sb[23:0];
  assign stage2_16_m0 = insn_o_1_680_0;
  assign insn_o_1_681_0 = stage2_16_pr[23:0];
  assign stage2_16_m1 = insn_o_1_681_0;
  assign insn_o_1_682_0 = stage2_16_sb[24:24];
  assign stage2_16_ms = insn_o_1_682_0;
  assign insn_o_1_683_0 = stage2_16_ms ? stage2_16_m1 : stage2_16_m0;
  assign stage2_16_mx = insn_o_1_683_0;
  assign insn_o_1_684_0 = stage2_zi_17[48:0];
  assign stage2_16_zl = insn_o_1_684_0;
  assign insn_o_1_685_0 = ~stage2_16_ms;
  assign stage2_16_zb = insn_o_1_685_0;
  assign insn_o_1_686_0 = {stage2_16_mx, stage2_16_zl, stage2_16_zb};
  assign insn_o_1_697_0 = stage2_zi_16[73:49];
  assign stage2_15_pr = insn_o_1_697_0;
  assign insn_o_1_698_0 = sub_663_d0;
  assign stage2_15_sb = insn_o_1_698_0;
  assign insn_o_1_699_0 = stage2_15_sb[23:0];
  assign stage2_15_m0 = insn_o_1_699_0;
  assign insn_o_1_700_0 = stage2_15_pr[23:0];
  assign stage2_15_m1 = insn_o_1_700_0;
  assign insn_o_1_701_0 = stage2_15_sb[24:24];
  assign stage2_15_ms = insn_o_1_701_0;
  assign insn_o_1_702_0 = stage2_15_ms ? stage2_15_m1 : stage2_15_m0;
  assign stage2_15_mx = insn_o_1_702_0;
  assign insn_o_1_703_0 = stage2_zi_16[48:0];
  assign stage2_15_zl = insn_o_1_703_0;
  assign insn_o_1_704_0 = ~stage2_15_ms;
  assign stage2_15_zb = insn_o_1_704_0;
  assign insn_o_1_705_0 = {stage2_15_mx, stage2_15_zl, stage2_15_zb};
  assign insn_o_1_716_0 = stage2_zi_15[73:49];
  assign stage2_14_pr = insn_o_1_716_0;
  assign insn_o_1_717_0 = sub_681_d0;
  assign stage2_14_sb = insn_o_1_717_0;
  assign insn_o_1_718_0 = stage2_14_sb[23:0];
  assign stage2_14_m0 = insn_o_1_718_0;
  assign insn_o_1_719_0 = stage2_14_pr[23:0];
  assign stage2_14_m1 = insn_o_1_719_0;
  assign insn_o_1_720_0 = stage2_14_sb[24:24];
  assign stage2_14_ms = insn_o_1_720_0;
  assign insn_o_1_721_0 = stage2_14_ms ? stage2_14_m1 : stage2_14_m0;
  assign stage2_14_mx = insn_o_1_721_0;
  assign insn_o_1_722_0 = stage2_zi_15[48:0];
  assign stage2_14_zl = insn_o_1_722_0;
  assign insn_o_1_723_0 = ~stage2_14_ms;
  assign stage2_14_zb = insn_o_1_723_0;
  assign insn_o_1_724_0 = {stage2_14_mx, stage2_14_zl, stage2_14_zb};
  assign insn_o_1_735_0 = stage2_zi_14[73:49];
  assign stage2_13_pr = insn_o_1_735_0;
  assign insn_o_1_736_0 = sub_699_d0;
  assign stage2_13_sb = insn_o_1_736_0;
  assign insn_o_1_737_0 = stage2_13_sb[23:0];
  assign stage2_13_m0 = insn_o_1_737_0;
  assign insn_o_1_738_0 = stage2_13_pr[23:0];
  assign stage2_13_m1 = insn_o_1_738_0;
  assign insn_o_1_739_0 = stage2_13_sb[24:24];
  assign stage2_13_ms = insn_o_1_739_0;
  assign insn_o_1_740_0 = stage2_13_ms ? stage2_13_m1 : stage2_13_m0;
  assign stage2_13_mx = insn_o_1_740_0;
  assign insn_o_1_741_0 = stage2_zi_14[48:0];
  assign stage2_13_zl = insn_o_1_741_0;
  assign insn_o_1_742_0 = ~stage2_13_ms;
  assign stage2_13_zb = insn_o_1_742_0;
  assign insn_o_1_743_0 = {stage2_13_mx, stage2_13_zl, stage2_13_zb};
  assign insn_o_1_754_0 = stage2_zi_13[73:49];
  assign stage2_12_pr = insn_o_1_754_0;
  assign insn_o_1_755_0 = sub_717_d0;
  assign stage2_12_sb = insn_o_1_755_0;
  assign insn_o_1_756_0 = stage2_12_sb[23:0];
  assign stage2_12_m0 = insn_o_1_756_0;
  assign insn_o_1_757_0 = stage2_12_pr[23:0];
  assign stage2_12_m1 = insn_o_1_757_0;
  assign insn_o_1_758_0 = stage2_12_sb[24:24];
  assign stage2_12_ms = insn_o_1_758_0;
  assign insn_o_1_759_0 = stage2_12_ms ? stage2_12_m1 : stage2_12_m0;
  assign stage2_12_mx = insn_o_1_759_0;
  assign insn_o_1_760_0 = stage2_zi_13[48:0];
  assign stage2_12_zl = insn_o_1_760_0;
  assign insn_o_1_761_0 = ~stage2_12_ms;
  assign stage2_12_zb = insn_o_1_761_0;
  assign insn_o_1_762_0 = {stage2_12_mx, stage2_12_zl, stage2_12_zb};
  assign insn_o_1_773_0 = stage2_zi_12[73:49];
  assign stage2_11_pr = insn_o_1_773_0;
  assign insn_o_1_774_0 = sub_735_d0;
  assign stage2_11_sb = insn_o_1_774_0;
  assign insn_o_1_775_0 = stage2_11_sb[23:0];
  assign stage2_11_m0 = insn_o_1_775_0;
  assign insn_o_1_776_0 = stage2_11_pr[23:0];
  assign stage2_11_m1 = insn_o_1_776_0;
  assign insn_o_1_777_0 = stage2_11_sb[24:24];
  assign stage2_11_ms = insn_o_1_777_0;
  assign insn_o_1_778_0 = stage2_11_ms ? stage2_11_m1 : stage2_11_m0;
  assign stage2_11_mx = insn_o_1_778_0;
  assign insn_o_1_779_0 = stage2_zi_12[48:0];
  assign stage2_11_zl = insn_o_1_779_0;
  assign insn_o_1_780_0 = ~stage2_11_ms;
  assign stage2_11_zb = insn_o_1_780_0;
  assign insn_o_1_781_0 = {stage2_11_mx, stage2_11_zl, stage2_11_zb};
  assign insn_o_1_792_0 = stage2_zi_11[73:49];
  assign stage2_10_pr = insn_o_1_792_0;
  assign insn_o_1_793_0 = sub_753_d0;
  assign stage2_10_sb = insn_o_1_793_0;
  assign insn_o_1_794_0 = stage2_10_sb[23:0];
  assign stage2_10_m0 = insn_o_1_794_0;
  assign insn_o_1_795_0 = stage2_10_pr[23:0];
  assign stage2_10_m1 = insn_o_1_795_0;
  assign insn_o_1_796_0 = stage2_10_sb[24:24];
  assign stage2_10_ms = insn_o_1_796_0;
  assign insn_o_1_797_0 = stage2_10_ms ? stage2_10_m1 : stage2_10_m0;
  assign stage2_10_mx = insn_o_1_797_0;
  assign insn_o_1_798_0 = stage2_zi_11[48:0];
  assign stage2_10_zl = insn_o_1_798_0;
  assign insn_o_1_799_0 = ~stage2_10_ms;
  assign stage2_10_zb = insn_o_1_799_0;
  assign insn_o_1_800_0 = {stage2_10_mx, stage2_10_zl, stage2_10_zb};
  assign insn_o_1_811_0 = stage2_zi_10[73:49];
  assign stage2_9_pr = insn_o_1_811_0;
  assign insn_o_1_812_0 = sub_771_d0;
  assign stage2_9_sb = insn_o_1_812_0;
  assign insn_o_1_813_0 = stage2_9_sb[23:0];
  assign stage2_9_m0 = insn_o_1_813_0;
  assign insn_o_1_814_0 = stage2_9_pr[23:0];
  assign stage2_9_m1 = insn_o_1_814_0;
  assign insn_o_1_815_0 = stage2_9_sb[24:24];
  assign stage2_9_ms = insn_o_1_815_0;
  assign insn_o_1_816_0 = stage2_9_ms ? stage2_9_m1 : stage2_9_m0;
  assign stage2_9_mx = insn_o_1_816_0;
  assign insn_o_1_817_0 = stage2_zi_10[48:0];
  assign stage2_9_zl = insn_o_1_817_0;
  assign insn_o_1_818_0 = ~stage2_9_ms;
  assign stage2_9_zb = insn_o_1_818_0;
  assign insn_o_1_819_0 = {stage2_9_mx, stage2_9_zl, stage2_9_zb};
  assign insn_o_1_830_0 = stage2_zi_09[73:49];
  assign stage2_8_pr = insn_o_1_830_0;
  assign insn_o_1_831_0 = sub_789_d0;
  assign stage2_8_sb = insn_o_1_831_0;
  assign insn_o_1_832_0 = stage2_8_sb[23:0];
  assign stage2_8_m0 = insn_o_1_832_0;
  assign insn_o_1_833_0 = stage2_8_pr[23:0];
  assign stage2_8_m1 = insn_o_1_833_0;
  assign insn_o_1_834_0 = stage2_8_sb[24:24];
  assign stage2_8_ms = insn_o_1_834_0;
  assign insn_o_1_835_0 = stage2_8_ms ? stage2_8_m1 : stage2_8_m0;
  assign stage2_8_mx = insn_o_1_835_0;
  assign insn_o_1_836_0 = stage2_zi_09[48:0];
  assign stage2_8_zl = insn_o_1_836_0;
  assign insn_o_1_837_0 = ~stage2_8_ms;
  assign stage2_8_zb = insn_o_1_837_0;
  assign insn_o_1_838_0 = {stage2_8_mx, stage2_8_zl, stage2_8_zb};
  assign insn_o_1_849_0 = stage2_zi_08[73:49];
  assign stage2_7_pr = insn_o_1_849_0;
  assign insn_o_1_850_0 = sub_807_d0;
  assign stage2_7_sb = insn_o_1_850_0;
  assign insn_o_1_851_0 = stage2_7_sb[23:0];
  assign stage2_7_m0 = insn_o_1_851_0;
  assign insn_o_1_852_0 = stage2_7_pr[23:0];
  assign stage2_7_m1 = insn_o_1_852_0;
  assign insn_o_1_853_0 = stage2_7_sb[24:24];
  assign stage2_7_ms = insn_o_1_853_0;
  assign insn_o_1_854_0 = stage2_7_ms ? stage2_7_m1 : stage2_7_m0;
  assign stage2_7_mx = insn_o_1_854_0;
  assign insn_o_1_855_0 = stage2_zi_08[48:0];
  assign stage2_7_zl = insn_o_1_855_0;
  assign insn_o_1_856_0 = ~stage2_7_ms;
  assign stage2_7_zb = insn_o_1_856_0;
  assign insn_o_1_857_0 = {stage2_7_mx, stage2_7_zl, stage2_7_zb};
  assign insn_o_1_868_0 = stage2_zi_07[73:49];
  assign stage2_6_pr = insn_o_1_868_0;
  assign insn_o_1_869_0 = sub_825_d0;
  assign stage2_6_sb = insn_o_1_869_0;
  assign insn_o_1_870_0 = stage2_6_sb[23:0];
  assign stage2_6_m0 = insn_o_1_870_0;
  assign insn_o_1_871_0 = stage2_6_pr[23:0];
  assign stage2_6_m1 = insn_o_1_871_0;
  assign insn_o_1_872_0 = stage2_6_sb[24:24];
  assign stage2_6_ms = insn_o_1_872_0;
  assign insn_o_1_873_0 = stage2_6_ms ? stage2_6_m1 : stage2_6_m0;
  assign stage2_6_mx = insn_o_1_873_0;
  assign insn_o_1_874_0 = stage2_zi_07[48:0];
  assign stage2_6_zl = insn_o_1_874_0;
  assign insn_o_1_875_0 = ~stage2_6_ms;
  assign stage2_6_zb = insn_o_1_875_0;
  assign insn_o_1_876_0 = {stage2_6_mx, stage2_6_zl, stage2_6_zb};
  assign insn_o_1_887_0 = stage2_zi_06[73:49];
  assign stage2_5_pr = insn_o_1_887_0;
  assign insn_o_1_888_0 = sub_843_d0;
  assign stage2_5_sb = insn_o_1_888_0;
  assign insn_o_1_889_0 = stage2_5_sb[23:0];
  assign stage2_5_m0 = insn_o_1_889_0;
  assign insn_o_1_890_0 = stage2_5_pr[23:0];
  assign stage2_5_m1 = insn_o_1_890_0;
  assign insn_o_1_891_0 = stage2_5_sb[24:24];
  assign stage2_5_ms = insn_o_1_891_0;
  assign insn_o_1_892_0 = stage2_5_ms ? stage2_5_m1 : stage2_5_m0;
  assign stage2_5_mx = insn_o_1_892_0;
  assign insn_o_1_893_0 = stage2_zi_06[48:0];
  assign stage2_5_zl = insn_o_1_893_0;
  assign insn_o_1_894_0 = ~stage2_5_ms;
  assign stage2_5_zb = insn_o_1_894_0;
  assign insn_o_1_895_0 = {stage2_5_mx, stage2_5_zl, stage2_5_zb};
  assign insn_o_1_906_0 = stage2_zi_05[73:49];
  assign stage2_4_pr = insn_o_1_906_0;
  assign insn_o_1_907_0 = sub_861_d0;
  assign stage2_4_sb = insn_o_1_907_0;
  assign insn_o_1_908_0 = stage2_4_sb[23:0];
  assign stage2_4_m0 = insn_o_1_908_0;
  assign insn_o_1_909_0 = stage2_4_pr[23:0];
  assign stage2_4_m1 = insn_o_1_909_0;
  assign insn_o_1_910_0 = stage2_4_sb[24:24];
  assign stage2_4_ms = insn_o_1_910_0;
  assign insn_o_1_911_0 = stage2_4_ms ? stage2_4_m1 : stage2_4_m0;
  assign stage2_4_mx = insn_o_1_911_0;
  assign insn_o_1_912_0 = stage2_zi_05[48:0];
  assign stage2_4_zl = insn_o_1_912_0;
  assign insn_o_1_913_0 = ~stage2_4_ms;
  assign stage2_4_zb = insn_o_1_913_0;
  assign insn_o_1_914_0 = {stage2_4_mx, stage2_4_zl, stage2_4_zb};
  assign insn_o_1_925_0 = stage2_zi_04[73:49];
  assign stage2_3_pr = insn_o_1_925_0;
  assign insn_o_1_926_0 = sub_879_d0;
  assign stage2_3_sb = insn_o_1_926_0;
  assign insn_o_1_927_0 = stage2_3_sb[23:0];
  assign stage2_3_m0 = insn_o_1_927_0;
  assign insn_o_1_928_0 = stage2_3_pr[23:0];
  assign stage2_3_m1 = insn_o_1_928_0;
  assign insn_o_1_929_0 = stage2_3_sb[24:24];
  assign stage2_3_ms = insn_o_1_929_0;
  assign insn_o_1_930_0 = stage2_3_ms ? stage2_3_m1 : stage2_3_m0;
  assign stage2_3_mx = insn_o_1_930_0;
  assign insn_o_1_931_0 = stage2_zi_04[48:0];
  assign stage2_3_zl = insn_o_1_931_0;
  assign insn_o_1_932_0 = ~stage2_3_ms;
  assign stage2_3_zb = insn_o_1_932_0;
  assign insn_o_1_933_0 = {stage2_3_mx, stage2_3_zl, stage2_3_zb};
  assign insn_o_1_944_0 = stage2_zi_03[73:49];
  assign stage2_2_pr = insn_o_1_944_0;
  assign insn_o_1_945_0 = sub_897_d0;
  assign stage2_2_sb = insn_o_1_945_0;
  assign insn_o_1_946_0 = stage2_2_sb[23:0];
  assign stage2_2_m0 = insn_o_1_946_0;
  assign insn_o_1_947_0 = stage2_2_pr[23:0];
  assign stage2_2_m1 = insn_o_1_947_0;
  assign insn_o_1_948_0 = stage2_2_sb[24:24];
  assign stage2_2_ms = insn_o_1_948_0;
  assign insn_o_1_949_0 = stage2_2_ms ? stage2_2_m1 : stage2_2_m0;
  assign stage2_2_mx = insn_o_1_949_0;
  assign insn_o_1_950_0 = stage2_zi_03[48:0];
  assign stage2_2_zl = insn_o_1_950_0;
  assign insn_o_1_951_0 = ~stage2_2_ms;
  assign stage2_2_zb = insn_o_1_951_0;
  assign insn_o_1_952_0 = {stage2_2_mx, stage2_2_zl, stage2_2_zb};
  assign insn_o_1_963_0 = stage2_zi_02[73:49];
  assign stage2_1_pr = insn_o_1_963_0;
  assign insn_o_1_964_0 = sub_915_d0;
  assign stage2_1_sb = insn_o_1_964_0;
  assign insn_o_1_965_0 = stage2_1_sb[23:0];
  assign stage2_1_m0 = insn_o_1_965_0;
  assign insn_o_1_966_0 = stage2_1_pr[23:0];
  assign stage2_1_m1 = insn_o_1_966_0;
  assign insn_o_1_967_0 = stage2_1_sb[24:24];
  assign stage2_1_ms = insn_o_1_967_0;
  assign insn_o_1_968_0 = stage2_1_ms ? stage2_1_m1 : stage2_1_m0;
  assign stage2_1_mx = insn_o_1_968_0;
  assign insn_o_1_969_0 = stage2_zi_02[48:0];
  assign stage2_1_zl = insn_o_1_969_0;
  assign insn_o_1_970_0 = ~stage2_1_ms;
  assign stage2_1_zb = insn_o_1_970_0;
  assign insn_o_1_971_0 = {stage2_1_mx, stage2_1_zl, stage2_1_zb};
  assign insn_o_1_982_0 = stage2_zi_01[73:49];
  assign stage2_0_pr = insn_o_1_982_0;
  assign insn_o_1_983_0 = sub_933_d0;
  assign stage2_0_sb = insn_o_1_983_0;
  assign insn_o_1_984_0 = stage2_0_sb[23:0];
  assign stage2_0_m0 = insn_o_1_984_0;
  assign insn_o_1_985_0 = stage2_0_pr[23:0];
  assign stage2_0_m1 = insn_o_1_985_0;
  assign insn_o_1_986_0 = stage2_0_sb[24:24];
  assign stage2_0_ms = insn_o_1_986_0;
  assign insn_o_1_987_0 = stage2_0_ms ? stage2_0_m1 : stage2_0_m0;
  assign stage2_0_mx = insn_o_1_987_0;
  assign insn_o_1_988_0 = stage2_zi_01[48:0];
  assign stage2_0_zl = insn_o_1_988_0;
  assign insn_o_1_989_0 = ~stage2_0_ms;
  assign stage2_0_zb = insn_o_1_989_0;
  assign insn_o_1_990_0 = {stage2_0_mx, stage2_0_zl, stage2_0_zb};
  assign insn_o_1_999_0 = add_949_d0;
  assign insn_o_1_1001_0 = stage2_zi_00[25:25];
  assign stage3_z_msb = insn_o_1_1001_0;
  assign insn_o_1_1002_0 = stage2_zi_00[24:0];
  assign anon_1008 = insn_o_1_1002_0;
  assign insn_o_1_1003_0 = {anon_1008, 2'd3};
  assign anon_1009 = insn_o_1_1003_0;
  assign insn_o_1_1004_0 = stage2_zi_00[25:0];
  assign anon_1010 = insn_o_1_1004_0;
  assign insn_o_1_1005_0 = {anon_1010, 1'd1};
  assign anon_1011 = insn_o_1_1005_0;
  assign insn_o_1_1006_0 = stage3_z_msb ? anon_1011 : anon_1009;
  assign insn_o_1_1007_0 = ~stage3_z_msb;
  assign anon_1012 = insn_o_1_1007_0;
  assign insn_o_1_1008_0 = sub_957_d0;
  assign insn_o_1_1016_0 = stage3_fraction[26:3];
  assign stage4_fraction_data = insn_o_1_1016_0;
  assign insn_o_1_1017_0 = stage3_fraction[3:3];
  assign stage4_s_least = insn_o_1_1017_0;
  assign insn_o_1_1018_0 = stage3_fraction[2:2];
  assign stage4_s_guard = insn_o_1_1018_0;
  assign insn_o_1_1019_0 = stage3_fraction[1:1];
  assign stage4_s_round = insn_o_1_1019_0;
  assign insn_o_1_1020_0 = stage3_fraction[0:0];
  assign stage4_s_sticky = insn_o_1_1020_0;
  assign insn_o_1_1021_0 = stage4_s_least | stage4_s_round;
  assign anon_1026 = insn_o_1_1021_0;
  assign insn_o_1_1022_0 = anon_1026 | stage4_s_sticky;
  assign anon_1027 = insn_o_1_1022_0;
  assign insn_o_1_1023_0 = stage4_s_guard & anon_1027;
  assign stage4_increment = insn_o_1_1023_0;
  assign insn_o_1_1024_0 = add_973_d0;
  assign insn_o_1_1025_0 = eq_974_d0;
  assign anon_1028 = insn_o_1_1025_0;
  assign insn_o_1_1026_0 = stage4_increment & anon_1028;
  assign anon_1029 = insn_o_1_1026_0;
  assign insn_o_1_1027_0 = add_976_d0;
  assign insn_o_1_1035_0 = gt_984_d0;
  assign stage5_exp_natural = insn_o_1_1035_0;
  assign insn_o_1_1036_0 = ~stage5_exp_natural;
  assign stage5_exp_underflow = insn_o_1_1036_0;
  assign insn_o_1_1037_0 = gte_986_d0;
  assign stage5_exp_overflow = insn_o_1_1037_0;
  assign insn_o_1_1038_0 = stage4_exponent[7:0];
  assign stage5_exponent_in = insn_o_1_1038_0;
  assign insn_o_1_1039_0 = stage4_fraction[22:0];
  assign stage5_fraction_in = insn_o_1_1039_0;
  assign insn_o_1_1040_0 = stage5_exp_overflow ? 8'd255 : stage5_exponent_in;
  assign stage5_exponent_i1 = insn_o_1_1040_0;
  assign insn_o_1_1041_0 = stage5_exp_overflow ? 23'd0 : stage5_fraction_in;
  assign stage5_fraction_i1 = insn_o_1_1041_0;
  assign insn_o_1_1042_0 = stage5_exp_underflow ? 8'd0 : stage5_exponent_i1;
  assign stage5_exponent_di = insn_o_1_1042_0;
  assign insn_o_1_1043_0 = stage5_exp_underflow ? 23'd0 : stage5_fraction_i1;
  assign stage5_fraction_di = insn_o_1_1043_0;
  assign stage5_a_is_zero = stage4_a_is_zero;
  assign stage5_a_is_inf = stage4_a_is_inf;
  assign stage5_a_is_nan = stage4_a_is_nan;
  assign insn_o_1_1047_0 = stage5_a_is_zero | stage5_a_is_inf;
  assign anon_1056 = insn_o_1_1047_0;
  assign insn_o_1_1048_0 = anon_1056 | stage5_a_is_nan;
  assign anon_1057 = insn_o_1_1048_0;
  assign insn_o_1_1049_0 = ~anon_1057;
  assign stage5_a_is_norm = insn_o_1_1049_0;
  assign stage5_b_is_zero = stage4_b_is_zero;
  assign stage5_b_is_inf = stage4_b_is_inf;
  assign stage5_b_is_nan = stage4_b_is_nan;
  assign insn_o_1_1053_0 = stage5_b_is_zero | stage5_b_is_inf;
  assign anon_1062 = insn_o_1_1053_0;
  assign insn_o_1_1054_0 = anon_1062 | stage5_b_is_nan;
  assign anon_1063 = insn_o_1_1054_0;
  assign insn_o_1_1055_0 = ~anon_1063;
  assign stage5_b_is_norm = insn_o_1_1055_0;
  assign insn_o_1_1056_0 = stage5_a_is_zero & stage5_b_is_inf;
  assign anon_1065 = insn_o_1_1056_0;
  assign insn_o_1_1057_0 = stage5_a_is_zero & stage5_b_is_norm;
  assign anon_1066 = insn_o_1_1057_0;
  assign insn_o_1_1058_0 = anon_1065 | anon_1066;
  assign anon_1067 = insn_o_1_1058_0;
  assign insn_o_1_1059_0 = stage5_a_is_norm & stage5_b_is_inf;
  assign anon_1068 = insn_o_1_1059_0;
  assign insn_o_1_1060_0 = anon_1067 | anon_1068;
  assign stage5_set_zero = insn_o_1_1060_0;
  assign insn_o_1_1061_0 = stage5_a_is_inf & stage5_b_is_zero;
  assign anon_1070 = insn_o_1_1061_0;
  assign insn_o_1_1062_0 = stage5_a_is_inf & stage5_b_is_norm;
  assign anon_1071 = insn_o_1_1062_0;
  assign insn_o_1_1063_0 = anon_1070 | anon_1071;
  assign anon_1072 = insn_o_1_1063_0;
  assign insn_o_1_1064_0 = stage5_a_is_norm & stage5_b_is_zero;
  assign anon_1073 = insn_o_1_1064_0;
  assign insn_o_1_1065_0 = anon_1072 | anon_1073;
  assign stage5_set_inf = insn_o_1_1065_0;
  assign insn_o_1_1066_0 = stage5_a_is_norm & stage5_b_is_norm;
  assign stage5_set_norm = insn_o_1_1066_0;
  assign insn_o_1_1067_0 = stage5_a_is_zero & stage5_b_is_zero;
  assign anon_1076 = insn_o_1_1067_0;
  assign insn_o_1_1068_0 = stage5_a_is_zero & stage5_b_is_nan;
  assign anon_1077 = insn_o_1_1068_0;
  assign insn_o_1_1069_0 = anon_1076 | anon_1077;
  assign anon_1078 = insn_o_1_1069_0;
  assign insn_o_1_1070_0 = stage5_a_is_inf & stage5_b_is_inf;
  assign anon_1079 = insn_o_1_1070_0;
  assign insn_o_1_1071_0 = anon_1078 | anon_1079;
  assign anon_1080 = insn_o_1_1071_0;
  assign insn_o_1_1072_0 = stage5_a_is_inf & stage5_b_is_nan;
  assign anon_1081 = insn_o_1_1072_0;
  assign insn_o_1_1073_0 = anon_1080 | anon_1081;
  assign anon_1082 = insn_o_1_1073_0;
  assign insn_o_1_1074_0 = anon_1082 | stage5_a_is_nan;
  assign anon_1083 = insn_o_1_1074_0;
  assign insn_o_1_1075_0 = stage5_a_is_norm & stage5_b_is_nan;
  assign anon_1084 = insn_o_1_1075_0;
  assign insn_o_1_1076_0 = anon_1083 | anon_1084;
  assign stage5_set_nan = insn_o_1_1076_0;
  assign insn_o_1_1077_0 = stage5_set_norm ? stage5_fraction_di : 23'd2097152;
  assign stage5_fraction_o0 = insn_o_1_1077_0;
  assign insn_o_1_1078_0 = stage5_set_norm ? stage5_exponent_di : 8'd255;
  assign stage5_exponent_o0 = insn_o_1_1078_0;
  assign insn_o_1_1079_0 = stage5_set_inf ? 23'd0 : stage5_fraction_o0;
  assign stage5_fraction_o1 = insn_o_1_1079_0;
  assign insn_o_1_1080_0 = stage5_set_inf ? 8'd255 : stage5_exponent_o0;
  assign stage5_exponent_o1 = insn_o_1_1080_0;
  assign insn_o_1_1081_0 = stage5_set_nan ? 1'd0 : stage4_sign;
  assign stage5_sign_o = insn_o_1_1081_0;
  assign insn_o_1_1082_0 = stage5_set_zero ? 23'd0 : stage5_fraction_o1;
  assign stage5_fraction_o = insn_o_1_1082_0;
  assign insn_o_1_1083_0 = stage5_set_zero ? 8'd0 : stage5_exponent_o1;
  assign stage5_exponent_o = insn_o_1_1083_0;
  assign insn_o_1_1084_0 = {stage5_sign_o, stage5_exponent_o, stage5_fraction_o};
  assign stage5_result = insn_o_1_1084_0;

  // Table 1
  always @(posedge clk) begin
    if (!rst_n) begin
      st_1_1 <= 0;
      st_1_2 <= 0;
      st_1_3 <= 0;
      st_1_4 <= 0;
      st_1_5 <= 0;
      st_1_6 <= 0;
      st_1_7 <= 0;
      st_1_8 <= 0;
      st_1_9 <= 0;
      st_1_10 <= 0;
      st_1_11 <= 0;
      st_1_12 <= 0;
      st_1_13 <= 0;
      st_1_14 <= 0;
      st_1_15 <= 0;
      st_1_16 <= 0;
      st_1_17 <= 0;
      st_1_18 <= 0;
      st_1_19 <= 0;
      st_1_20 <= 0;
      st_1_21 <= 0;
      st_1_22 <= 0;
      st_1_23 <= 0;
      st_1_24 <= 0;
      st_1_25 <= 0;
      st_1_26 <= 0;
      st_1_27 <= 0;
      st_1_28 <= 0;
      st_1_29 <= 0;
      st_1_30 <= 0;
      st_1_31 <= 0;
      st_1_32 <= 0;
      st_1_33 <= 0;
      st_1_34 <= 0;
      st_1_35 <= 0;
      st_1_36 <= 0;
      st_1_37 <= 0;
      st_1_38 <= 0;
      st_1_39 <= 0;
      st_1_40 <= 0;
      st_1_41 <= 0;
      st_1_42 <= 0;
      st_1_43 <= 0;
      st_1_44 <= 0;
      st_1_45 <= 0;
      st_1_46 <= 0;
      st_1_47 <= 0;
      st_1_48 <= 0;
      st_1_49 <= 0;
      st_1_50 <= 0;
      st_1_51 <= 0;
      st_1_52 <= 0;
      st_1_53 <= 0;
      st_1_54 <= 0;
      st_1_55 <= 0;
    end else begin
      z_valid <= ((st_1_55) ? 1'd1 : 0);
      if (start) begin
          stage1_a_exponent <= stage1_a_exponent_in;
          stage1_a_sign <= stage1_a_sign_in;
          stage1_a_exponent_is_all_0 <= stage1_a_exponent_zero;
          stage1_b_exponent <= stage1_b_exponent_in;
          stage1_b_sign <= stage1_b_sign_in;
          stage1_b_exponent_is_all_0 <= stage1_b_exponent_zero;
          stage1_a_fraction <= insn_o_1_11_0;
          stage1_a_fraction_is_all_0 <= insn_o_1_15_0;
          stage1_b_fraction <= insn_o_1_22_0;
          stage1_b_fraction_is_all_0 <= insn_o_1_26_0;
      end
      st_1_2 <= start;
      if (st_1_2) begin
          stage2_di_50 <= stage1_b_fraction;
          stage2_zi_50 <= insn_o_1_32_0;
          stage2_exponent_50 <= insn_o_1_34_0;
          stage2_sign_50 <= insn_o_1_35_0;
          stage2_a_is_zero_50 <= insn_o_1_40_0;
          stage2_a_is_inf_50 <= insn_o_1_41_0;
          stage2_a_is_nan_50 <= insn_o_1_42_0;
          stage2_b_is_zero_50 <= insn_o_1_47_0;
          stage2_b_is_inf_50 <= insn_o_1_48_0;
          stage2_b_is_nan_50 <= insn_o_1_49_0;
      end
      st_1_3 <= st_1_2;
      if (st_1_3) begin
          stage2_di_49 <= stage2_di_50;
          stage2_sign_49 <= stage2_sign_50;
          stage2_a_is_zero_49 <= stage2_a_is_zero_50;
          stage2_a_is_inf_49 <= stage2_a_is_inf_50;
          stage2_a_is_nan_49 <= stage2_a_is_nan_50;
          stage2_b_is_zero_49 <= stage2_b_is_zero_50;
          stage2_b_is_inf_49 <= stage2_b_is_inf_50;
          stage2_b_is_nan_49 <= stage2_b_is_nan_50;
          stage2_exponent_49 <= stage2_exponent_50;
          stage2_zi_49 <= insn_o_1_59_0;
      end
      st_1_4 <= st_1_3;
      if (st_1_4) begin
          stage2_di_48 <= stage2_di_49;
          stage2_sign_48 <= stage2_sign_49;
          stage2_a_is_zero_48 <= stage2_a_is_zero_49;
          stage2_a_is_inf_48 <= stage2_a_is_inf_49;
          stage2_a_is_nan_48 <= stage2_a_is_nan_49;
          stage2_b_is_zero_48 <= stage2_b_is_zero_49;
          stage2_b_is_inf_48 <= stage2_b_is_inf_49;
          stage2_b_is_nan_48 <= stage2_b_is_nan_49;
          stage2_exponent_48 <= stage2_exponent_49;
          stage2_zi_48 <= insn_o_1_78_0;
      end
      st_1_5 <= st_1_4;
      if (st_1_5) begin
          stage2_di_47 <= stage2_di_48;
          stage2_sign_47 <= stage2_sign_48;
          stage2_a_is_zero_47 <= stage2_a_is_zero_48;
          stage2_a_is_inf_47 <= stage2_a_is_inf_48;
          stage2_a_is_nan_47 <= stage2_a_is_nan_48;
          stage2_b_is_zero_47 <= stage2_b_is_zero_48;
          stage2_b_is_inf_47 <= stage2_b_is_inf_48;
          stage2_b_is_nan_47 <= stage2_b_is_nan_48;
          stage2_exponent_47 <= stage2_exponent_48;
          stage2_zi_47 <= insn_o_1_97_0;
      end
      st_1_6 <= st_1_5;
      if (st_1_6) begin
          stage2_di_46 <= stage2_di_47;
          stage2_sign_46 <= stage2_sign_47;
          stage2_a_is_zero_46 <= stage2_a_is_zero_47;
          stage2_a_is_inf_46 <= stage2_a_is_inf_47;
          stage2_a_is_nan_46 <= stage2_a_is_nan_47;
          stage2_b_is_zero_46 <= stage2_b_is_zero_47;
          stage2_b_is_inf_46 <= stage2_b_is_inf_47;
          stage2_b_is_nan_46 <= stage2_b_is_nan_47;
          stage2_exponent_46 <= stage2_exponent_47;
          stage2_zi_46 <= insn_o_1_116_0;
      end
      st_1_7 <= st_1_6;
      if (st_1_7) begin
          stage2_di_45 <= stage2_di_46;
          stage2_sign_45 <= stage2_sign_46;
          stage2_a_is_zero_45 <= stage2_a_is_zero_46;
          stage2_a_is_inf_45 <= stage2_a_is_inf_46;
          stage2_a_is_nan_45 <= stage2_a_is_nan_46;
          stage2_b_is_zero_45 <= stage2_b_is_zero_46;
          stage2_b_is_inf_45 <= stage2_b_is_inf_46;
          stage2_b_is_nan_45 <= stage2_b_is_nan_46;
          stage2_exponent_45 <= stage2_exponent_46;
          stage2_zi_45 <= insn_o_1_135_0;
      end
      st_1_8 <= st_1_7;
      if (st_1_8) begin
          stage2_di_44 <= stage2_di_45;
          stage2_sign_44 <= stage2_sign_45;
          stage2_a_is_zero_44 <= stage2_a_is_zero_45;
          stage2_a_is_inf_44 <= stage2_a_is_inf_45;
          stage2_a_is_nan_44 <= stage2_a_is_nan_45;
          stage2_b_is_zero_44 <= stage2_b_is_zero_45;
          stage2_b_is_inf_44 <= stage2_b_is_inf_45;
          stage2_b_is_nan_44 <= stage2_b_is_nan_45;
          stage2_exponent_44 <= stage2_exponent_45;
          stage2_zi_44 <= insn_o_1_154_0;
      end
      st_1_9 <= st_1_8;
      if (st_1_9) begin
          stage2_di_43 <= stage2_di_44;
          stage2_sign_43 <= stage2_sign_44;
          stage2_a_is_zero_43 <= stage2_a_is_zero_44;
          stage2_a_is_inf_43 <= stage2_a_is_inf_44;
          stage2_a_is_nan_43 <= stage2_a_is_nan_44;
          stage2_b_is_zero_43 <= stage2_b_is_zero_44;
          stage2_b_is_inf_43 <= stage2_b_is_inf_44;
          stage2_b_is_nan_43 <= stage2_b_is_nan_44;
          stage2_exponent_43 <= stage2_exponent_44;
          stage2_zi_43 <= insn_o_1_173_0;
      end
      st_1_10 <= st_1_9;
      if (st_1_10) begin
          stage2_di_42 <= stage2_di_43;
          stage2_sign_42 <= stage2_sign_43;
          stage2_a_is_zero_42 <= stage2_a_is_zero_43;
          stage2_a_is_inf_42 <= stage2_a_is_inf_43;
          stage2_a_is_nan_42 <= stage2_a_is_nan_43;
          stage2_b_is_zero_42 <= stage2_b_is_zero_43;
          stage2_b_is_inf_42 <= stage2_b_is_inf_43;
          stage2_b_is_nan_42 <= stage2_b_is_nan_43;
          stage2_exponent_42 <= stage2_exponent_43;
          stage2_zi_42 <= insn_o_1_192_0;
      end
      st_1_11 <= st_1_10;
      if (st_1_11) begin
          stage2_di_41 <= stage2_di_42;
          stage2_sign_41 <= stage2_sign_42;
          stage2_a_is_zero_41 <= stage2_a_is_zero_42;
          stage2_a_is_inf_41 <= stage2_a_is_inf_42;
          stage2_a_is_nan_41 <= stage2_a_is_nan_42;
          stage2_b_is_zero_41 <= stage2_b_is_zero_42;
          stage2_b_is_inf_41 <= stage2_b_is_inf_42;
          stage2_b_is_nan_41 <= stage2_b_is_nan_42;
          stage2_exponent_41 <= stage2_exponent_42;
          stage2_zi_41 <= insn_o_1_211_0;
      end
      st_1_12 <= st_1_11;
      if (st_1_12) begin
          stage2_di_40 <= stage2_di_41;
          stage2_sign_40 <= stage2_sign_41;
          stage2_a_is_zero_40 <= stage2_a_is_zero_41;
          stage2_a_is_inf_40 <= stage2_a_is_inf_41;
          stage2_a_is_nan_40 <= stage2_a_is_nan_41;
          stage2_b_is_zero_40 <= stage2_b_is_zero_41;
          stage2_b_is_inf_40 <= stage2_b_is_inf_41;
          stage2_b_is_nan_40 <= stage2_b_is_nan_41;
          stage2_exponent_40 <= stage2_exponent_41;
          stage2_zi_40 <= insn_o_1_230_0;
      end
      st_1_13 <= st_1_12;
      if (st_1_13) begin
          stage2_di_39 <= stage2_di_40;
          stage2_sign_39 <= stage2_sign_40;
          stage2_a_is_zero_39 <= stage2_a_is_zero_40;
          stage2_a_is_inf_39 <= stage2_a_is_inf_40;
          stage2_a_is_nan_39 <= stage2_a_is_nan_40;
          stage2_b_is_zero_39 <= stage2_b_is_zero_40;
          stage2_b_is_inf_39 <= stage2_b_is_inf_40;
          stage2_b_is_nan_39 <= stage2_b_is_nan_40;
          stage2_exponent_39 <= stage2_exponent_40;
          stage2_zi_39 <= insn_o_1_249_0;
      end
      st_1_14 <= st_1_13;
      if (st_1_14) begin
          stage2_di_38 <= stage2_di_39;
          stage2_sign_38 <= stage2_sign_39;
          stage2_a_is_zero_38 <= stage2_a_is_zero_39;
          stage2_a_is_inf_38 <= stage2_a_is_inf_39;
          stage2_a_is_nan_38 <= stage2_a_is_nan_39;
          stage2_b_is_zero_38 <= stage2_b_is_zero_39;
          stage2_b_is_inf_38 <= stage2_b_is_inf_39;
          stage2_b_is_nan_38 <= stage2_b_is_nan_39;
          stage2_exponent_38 <= stage2_exponent_39;
          stage2_zi_38 <= insn_o_1_268_0;
      end
      st_1_15 <= st_1_14;
      if (st_1_15) begin
          stage2_di_37 <= stage2_di_38;
          stage2_sign_37 <= stage2_sign_38;
          stage2_a_is_zero_37 <= stage2_a_is_zero_38;
          stage2_a_is_inf_37 <= stage2_a_is_inf_38;
          stage2_a_is_nan_37 <= stage2_a_is_nan_38;
          stage2_b_is_zero_37 <= stage2_b_is_zero_38;
          stage2_b_is_inf_37 <= stage2_b_is_inf_38;
          stage2_b_is_nan_37 <= stage2_b_is_nan_38;
          stage2_exponent_37 <= stage2_exponent_38;
          stage2_zi_37 <= insn_o_1_287_0;
      end
      st_1_16 <= st_1_15;
      if (st_1_16) begin
          stage2_di_36 <= stage2_di_37;
          stage2_sign_36 <= stage2_sign_37;
          stage2_a_is_zero_36 <= stage2_a_is_zero_37;
          stage2_a_is_inf_36 <= stage2_a_is_inf_37;
          stage2_a_is_nan_36 <= stage2_a_is_nan_37;
          stage2_b_is_zero_36 <= stage2_b_is_zero_37;
          stage2_b_is_inf_36 <= stage2_b_is_inf_37;
          stage2_b_is_nan_36 <= stage2_b_is_nan_37;
          stage2_exponent_36 <= stage2_exponent_37;
          stage2_zi_36 <= insn_o_1_306_0;
      end
      st_1_17 <= st_1_16;
      if (st_1_17) begin
          stage2_di_35 <= stage2_di_36;
          stage2_sign_35 <= stage2_sign_36;
          stage2_a_is_zero_35 <= stage2_a_is_zero_36;
          stage2_a_is_inf_35 <= stage2_a_is_inf_36;
          stage2_a_is_nan_35 <= stage2_a_is_nan_36;
          stage2_b_is_zero_35 <= stage2_b_is_zero_36;
          stage2_b_is_inf_35 <= stage2_b_is_inf_36;
          stage2_b_is_nan_35 <= stage2_b_is_nan_36;
          stage2_exponent_35 <= stage2_exponent_36;
          stage2_zi_35 <= insn_o_1_325_0;
      end
      st_1_18 <= st_1_17;
      if (st_1_18) begin
          stage2_di_34 <= stage2_di_35;
          stage2_sign_34 <= stage2_sign_35;
          stage2_a_is_zero_34 <= stage2_a_is_zero_35;
          stage2_a_is_inf_34 <= stage2_a_is_inf_35;
          stage2_a_is_nan_34 <= stage2_a_is_nan_35;
          stage2_b_is_zero_34 <= stage2_b_is_zero_35;
          stage2_b_is_inf_34 <= stage2_b_is_inf_35;
          stage2_b_is_nan_34 <= stage2_b_is_nan_35;
          stage2_exponent_34 <= stage2_exponent_35;
          stage2_zi_34 <= insn_o_1_344_0;
      end
      st_1_19 <= st_1_18;
      if (st_1_19) begin
          stage2_di_33 <= stage2_di_34;
          stage2_sign_33 <= stage2_sign_34;
          stage2_a_is_zero_33 <= stage2_a_is_zero_34;
          stage2_a_is_inf_33 <= stage2_a_is_inf_34;
          stage2_a_is_nan_33 <= stage2_a_is_nan_34;
          stage2_b_is_zero_33 <= stage2_b_is_zero_34;
          stage2_b_is_inf_33 <= stage2_b_is_inf_34;
          stage2_b_is_nan_33 <= stage2_b_is_nan_34;
          stage2_exponent_33 <= stage2_exponent_34;
          stage2_zi_33 <= insn_o_1_363_0;
      end
      st_1_20 <= st_1_19;
      if (st_1_20) begin
          stage2_di_32 <= stage2_di_33;
          stage2_sign_32 <= stage2_sign_33;
          stage2_a_is_zero_32 <= stage2_a_is_zero_33;
          stage2_a_is_inf_32 <= stage2_a_is_inf_33;
          stage2_a_is_nan_32 <= stage2_a_is_nan_33;
          stage2_b_is_zero_32 <= stage2_b_is_zero_33;
          stage2_b_is_inf_32 <= stage2_b_is_inf_33;
          stage2_b_is_nan_32 <= stage2_b_is_nan_33;
          stage2_exponent_32 <= stage2_exponent_33;
          stage2_zi_32 <= insn_o_1_382_0;
      end
      st_1_21 <= st_1_20;
      if (st_1_21) begin
          stage2_di_31 <= stage2_di_32;
          stage2_sign_31 <= stage2_sign_32;
          stage2_a_is_zero_31 <= stage2_a_is_zero_32;
          stage2_a_is_inf_31 <= stage2_a_is_inf_32;
          stage2_a_is_nan_31 <= stage2_a_is_nan_32;
          stage2_b_is_zero_31 <= stage2_b_is_zero_32;
          stage2_b_is_inf_31 <= stage2_b_is_inf_32;
          stage2_b_is_nan_31 <= stage2_b_is_nan_32;
          stage2_exponent_31 <= stage2_exponent_32;
          stage2_zi_31 <= insn_o_1_401_0;
      end
      st_1_22 <= st_1_21;
      if (st_1_22) begin
          stage2_di_30 <= stage2_di_31;
          stage2_sign_30 <= stage2_sign_31;
          stage2_a_is_zero_30 <= stage2_a_is_zero_31;
          stage2_a_is_inf_30 <= stage2_a_is_inf_31;
          stage2_a_is_nan_30 <= stage2_a_is_nan_31;
          stage2_b_is_zero_30 <= stage2_b_is_zero_31;
          stage2_b_is_inf_30 <= stage2_b_is_inf_31;
          stage2_b_is_nan_30 <= stage2_b_is_nan_31;
          stage2_exponent_30 <= stage2_exponent_31;
          stage2_zi_30 <= insn_o_1_420_0;
      end
      st_1_23 <= st_1_22;
      if (st_1_23) begin
          stage2_di_29 <= stage2_di_30;
          stage2_sign_29 <= stage2_sign_30;
          stage2_a_is_zero_29 <= stage2_a_is_zero_30;
          stage2_a_is_inf_29 <= stage2_a_is_inf_30;
          stage2_a_is_nan_29 <= stage2_a_is_nan_30;
          stage2_b_is_zero_29 <= stage2_b_is_zero_30;
          stage2_b_is_inf_29 <= stage2_b_is_inf_30;
          stage2_b_is_nan_29 <= stage2_b_is_nan_30;
          stage2_exponent_29 <= stage2_exponent_30;
          stage2_zi_29 <= insn_o_1_439_0;
      end
      st_1_24 <= st_1_23;
      if (st_1_24) begin
          stage2_di_28 <= stage2_di_29;
          stage2_sign_28 <= stage2_sign_29;
          stage2_a_is_zero_28 <= stage2_a_is_zero_29;
          stage2_a_is_inf_28 <= stage2_a_is_inf_29;
          stage2_a_is_nan_28 <= stage2_a_is_nan_29;
          stage2_b_is_zero_28 <= stage2_b_is_zero_29;
          stage2_b_is_inf_28 <= stage2_b_is_inf_29;
          stage2_b_is_nan_28 <= stage2_b_is_nan_29;
          stage2_exponent_28 <= stage2_exponent_29;
          stage2_zi_28 <= insn_o_1_458_0;
      end
      st_1_25 <= st_1_24;
      if (st_1_25) begin
          stage2_di_27 <= stage2_di_28;
          stage2_sign_27 <= stage2_sign_28;
          stage2_a_is_zero_27 <= stage2_a_is_zero_28;
          stage2_a_is_inf_27 <= stage2_a_is_inf_28;
          stage2_a_is_nan_27 <= stage2_a_is_nan_28;
          stage2_b_is_zero_27 <= stage2_b_is_zero_28;
          stage2_b_is_inf_27 <= stage2_b_is_inf_28;
          stage2_b_is_nan_27 <= stage2_b_is_nan_28;
          stage2_exponent_27 <= stage2_exponent_28;
          stage2_zi_27 <= insn_o_1_477_0;
      end
      st_1_26 <= st_1_25;
      if (st_1_26) begin
          stage2_di_26 <= stage2_di_27;
          stage2_sign_26 <= stage2_sign_27;
          stage2_a_is_zero_26 <= stage2_a_is_zero_27;
          stage2_a_is_inf_26 <= stage2_a_is_inf_27;
          stage2_a_is_nan_26 <= stage2_a_is_nan_27;
          stage2_b_is_zero_26 <= stage2_b_is_zero_27;
          stage2_b_is_inf_26 <= stage2_b_is_inf_27;
          stage2_b_is_nan_26 <= stage2_b_is_nan_27;
          stage2_exponent_26 <= stage2_exponent_27;
          stage2_zi_26 <= insn_o_1_496_0;
      end
      st_1_27 <= st_1_26;
      if (st_1_27) begin
          stage2_di_25 <= stage2_di_26;
          stage2_sign_25 <= stage2_sign_26;
          stage2_a_is_zero_25 <= stage2_a_is_zero_26;
          stage2_a_is_inf_25 <= stage2_a_is_inf_26;
          stage2_a_is_nan_25 <= stage2_a_is_nan_26;
          stage2_b_is_zero_25 <= stage2_b_is_zero_26;
          stage2_b_is_inf_25 <= stage2_b_is_inf_26;
          stage2_b_is_nan_25 <= stage2_b_is_nan_26;
          stage2_exponent_25 <= stage2_exponent_26;
          stage2_zi_25 <= insn_o_1_515_0;
      end
      st_1_28 <= st_1_27;
      if (st_1_28) begin
          stage2_di_24 <= stage2_di_25;
          stage2_sign_24 <= stage2_sign_25;
          stage2_a_is_zero_24 <= stage2_a_is_zero_25;
          stage2_a_is_inf_24 <= stage2_a_is_inf_25;
          stage2_a_is_nan_24 <= stage2_a_is_nan_25;
          stage2_b_is_zero_24 <= stage2_b_is_zero_25;
          stage2_b_is_inf_24 <= stage2_b_is_inf_25;
          stage2_b_is_nan_24 <= stage2_b_is_nan_25;
          stage2_exponent_24 <= stage2_exponent_25;
          stage2_zi_24 <= insn_o_1_534_0;
      end
      st_1_29 <= st_1_28;
      if (st_1_29) begin
          stage2_di_23 <= stage2_di_24;
          stage2_sign_23 <= stage2_sign_24;
          stage2_a_is_zero_23 <= stage2_a_is_zero_24;
          stage2_a_is_inf_23 <= stage2_a_is_inf_24;
          stage2_a_is_nan_23 <= stage2_a_is_nan_24;
          stage2_b_is_zero_23 <= stage2_b_is_zero_24;
          stage2_b_is_inf_23 <= stage2_b_is_inf_24;
          stage2_b_is_nan_23 <= stage2_b_is_nan_24;
          stage2_exponent_23 <= stage2_exponent_24;
          stage2_zi_23 <= insn_o_1_553_0;
      end
      st_1_30 <= st_1_29;
      if (st_1_30) begin
          stage2_di_22 <= stage2_di_23;
          stage2_sign_22 <= stage2_sign_23;
          stage2_a_is_zero_22 <= stage2_a_is_zero_23;
          stage2_a_is_inf_22 <= stage2_a_is_inf_23;
          stage2_a_is_nan_22 <= stage2_a_is_nan_23;
          stage2_b_is_zero_22 <= stage2_b_is_zero_23;
          stage2_b_is_inf_22 <= stage2_b_is_inf_23;
          stage2_b_is_nan_22 <= stage2_b_is_nan_23;
          stage2_exponent_22 <= stage2_exponent_23;
          stage2_zi_22 <= insn_o_1_572_0;
      end
      st_1_31 <= st_1_30;
      if (st_1_31) begin
          stage2_di_21 <= stage2_di_22;
          stage2_sign_21 <= stage2_sign_22;
          stage2_a_is_zero_21 <= stage2_a_is_zero_22;
          stage2_a_is_inf_21 <= stage2_a_is_inf_22;
          stage2_a_is_nan_21 <= stage2_a_is_nan_22;
          stage2_b_is_zero_21 <= stage2_b_is_zero_22;
          stage2_b_is_inf_21 <= stage2_b_is_inf_22;
          stage2_b_is_nan_21 <= stage2_b_is_nan_22;
          stage2_exponent_21 <= stage2_exponent_22;
          stage2_zi_21 <= insn_o_1_591_0;
      end
      st_1_32 <= st_1_31;
      if (st_1_32) begin
          stage2_di_20 <= stage2_di_21;
          stage2_sign_20 <= stage2_sign_21;
          stage2_a_is_zero_20 <= stage2_a_is_zero_21;
          stage2_a_is_inf_20 <= stage2_a_is_inf_21;
          stage2_a_is_nan_20 <= stage2_a_is_nan_21;
          stage2_b_is_zero_20 <= stage2_b_is_zero_21;
          stage2_b_is_inf_20 <= stage2_b_is_inf_21;
          stage2_b_is_nan_20 <= stage2_b_is_nan_21;
          stage2_exponent_20 <= stage2_exponent_21;
          stage2_zi_20 <= insn_o_1_610_0;
      end
      st_1_33 <= st_1_32;
      if (st_1_33) begin
          stage2_di_19 <= stage2_di_20;
          stage2_sign_19 <= stage2_sign_20;
          stage2_a_is_zero_19 <= stage2_a_is_zero_20;
          stage2_a_is_inf_19 <= stage2_a_is_inf_20;
          stage2_a_is_nan_19 <= stage2_a_is_nan_20;
          stage2_b_is_zero_19 <= stage2_b_is_zero_20;
          stage2_b_is_inf_19 <= stage2_b_is_inf_20;
          stage2_b_is_nan_19 <= stage2_b_is_nan_20;
          stage2_exponent_19 <= stage2_exponent_20;
          stage2_zi_19 <= insn_o_1_629_0;
      end
      st_1_34 <= st_1_33;
      if (st_1_34) begin
          stage2_di_18 <= stage2_di_19;
          stage2_sign_18 <= stage2_sign_19;
          stage2_a_is_zero_18 <= stage2_a_is_zero_19;
          stage2_a_is_inf_18 <= stage2_a_is_inf_19;
          stage2_a_is_nan_18 <= stage2_a_is_nan_19;
          stage2_b_is_zero_18 <= stage2_b_is_zero_19;
          stage2_b_is_inf_18 <= stage2_b_is_inf_19;
          stage2_b_is_nan_18 <= stage2_b_is_nan_19;
          stage2_exponent_18 <= stage2_exponent_19;
          stage2_zi_18 <= insn_o_1_648_0;
      end
      st_1_35 <= st_1_34;
      if (st_1_35) begin
          stage2_di_17 <= stage2_di_18;
          stage2_sign_17 <= stage2_sign_18;
          stage2_a_is_zero_17 <= stage2_a_is_zero_18;
          stage2_a_is_inf_17 <= stage2_a_is_inf_18;
          stage2_a_is_nan_17 <= stage2_a_is_nan_18;
          stage2_b_is_zero_17 <= stage2_b_is_zero_18;
          stage2_b_is_inf_17 <= stage2_b_is_inf_18;
          stage2_b_is_nan_17 <= stage2_b_is_nan_18;
          stage2_exponent_17 <= stage2_exponent_18;
          stage2_zi_17 <= insn_o_1_667_0;
      end
      st_1_36 <= st_1_35;
      if (st_1_36) begin
          stage2_di_16 <= stage2_di_17;
          stage2_sign_16 <= stage2_sign_17;
          stage2_a_is_zero_16 <= stage2_a_is_zero_17;
          stage2_a_is_inf_16 <= stage2_a_is_inf_17;
          stage2_a_is_nan_16 <= stage2_a_is_nan_17;
          stage2_b_is_zero_16 <= stage2_b_is_zero_17;
          stage2_b_is_inf_16 <= stage2_b_is_inf_17;
          stage2_b_is_nan_16 <= stage2_b_is_nan_17;
          stage2_exponent_16 <= stage2_exponent_17;
          stage2_zi_16 <= insn_o_1_686_0;
      end
      st_1_37 <= st_1_36;
      if (st_1_37) begin
          stage2_di_15 <= stage2_di_16;
          stage2_sign_15 <= stage2_sign_16;
          stage2_a_is_zero_15 <= stage2_a_is_zero_16;
          stage2_a_is_inf_15 <= stage2_a_is_inf_16;
          stage2_a_is_nan_15 <= stage2_a_is_nan_16;
          stage2_b_is_zero_15 <= stage2_b_is_zero_16;
          stage2_b_is_inf_15 <= stage2_b_is_inf_16;
          stage2_b_is_nan_15 <= stage2_b_is_nan_16;
          stage2_exponent_15 <= stage2_exponent_16;
          stage2_zi_15 <= insn_o_1_705_0;
      end
      st_1_38 <= st_1_37;
      if (st_1_38) begin
          stage2_di_14 <= stage2_di_15;
          stage2_sign_14 <= stage2_sign_15;
          stage2_a_is_zero_14 <= stage2_a_is_zero_15;
          stage2_a_is_inf_14 <= stage2_a_is_inf_15;
          stage2_a_is_nan_14 <= stage2_a_is_nan_15;
          stage2_b_is_zero_14 <= stage2_b_is_zero_15;
          stage2_b_is_inf_14 <= stage2_b_is_inf_15;
          stage2_b_is_nan_14 <= stage2_b_is_nan_15;
          stage2_exponent_14 <= stage2_exponent_15;
          stage2_zi_14 <= insn_o_1_724_0;
      end
      st_1_39 <= st_1_38;
      if (st_1_39) begin
          stage2_di_13 <= stage2_di_14;
          stage2_sign_13 <= stage2_sign_14;
          stage2_a_is_zero_13 <= stage2_a_is_zero_14;
          stage2_a_is_inf_13 <= stage2_a_is_inf_14;
          stage2_a_is_nan_13 <= stage2_a_is_nan_14;
          stage2_b_is_zero_13 <= stage2_b_is_zero_14;
          stage2_b_is_inf_13 <= stage2_b_is_inf_14;
          stage2_b_is_nan_13 <= stage2_b_is_nan_14;
          stage2_exponent_13 <= stage2_exponent_14;
          stage2_zi_13 <= insn_o_1_743_0;
      end
      st_1_40 <= st_1_39;
      if (st_1_40) begin
          stage2_di_12 <= stage2_di_13;
          stage2_sign_12 <= stage2_sign_13;
          stage2_a_is_zero_12 <= stage2_a_is_zero_13;
          stage2_a_is_inf_12 <= stage2_a_is_inf_13;
          stage2_a_is_nan_12 <= stage2_a_is_nan_13;
          stage2_b_is_zero_12 <= stage2_b_is_zero_13;
          stage2_b_is_inf_12 <= stage2_b_is_inf_13;
          stage2_b_is_nan_12 <= stage2_b_is_nan_13;
          stage2_exponent_12 <= stage2_exponent_13;
          stage2_zi_12 <= insn_o_1_762_0;
      end
      st_1_41 <= st_1_40;
      if (st_1_41) begin
          stage2_di_11 <= stage2_di_12;
          stage2_sign_11 <= stage2_sign_12;
          stage2_a_is_zero_11 <= stage2_a_is_zero_12;
          stage2_a_is_inf_11 <= stage2_a_is_inf_12;
          stage2_a_is_nan_11 <= stage2_a_is_nan_12;
          stage2_b_is_zero_11 <= stage2_b_is_zero_12;
          stage2_b_is_inf_11 <= stage2_b_is_inf_12;
          stage2_b_is_nan_11 <= stage2_b_is_nan_12;
          stage2_exponent_11 <= stage2_exponent_12;
          stage2_zi_11 <= insn_o_1_781_0;
      end
      st_1_42 <= st_1_41;
      if (st_1_42) begin
          stage2_di_10 <= stage2_di_11;
          stage2_sign_10 <= stage2_sign_11;
          stage2_a_is_zero_10 <= stage2_a_is_zero_11;
          stage2_a_is_inf_10 <= stage2_a_is_inf_11;
          stage2_a_is_nan_10 <= stage2_a_is_nan_11;
          stage2_b_is_zero_10 <= stage2_b_is_zero_11;
          stage2_b_is_inf_10 <= stage2_b_is_inf_11;
          stage2_b_is_nan_10 <= stage2_b_is_nan_11;
          stage2_exponent_10 <= stage2_exponent_11;
          stage2_zi_10 <= insn_o_1_800_0;
      end
      st_1_43 <= st_1_42;
      if (st_1_43) begin
          stage2_di_09 <= stage2_di_10;
          stage2_sign_09 <= stage2_sign_10;
          stage2_a_is_zero_09 <= stage2_a_is_zero_10;
          stage2_a_is_inf_09 <= stage2_a_is_inf_10;
          stage2_a_is_nan_09 <= stage2_a_is_nan_10;
          stage2_b_is_zero_09 <= stage2_b_is_zero_10;
          stage2_b_is_inf_09 <= stage2_b_is_inf_10;
          stage2_b_is_nan_09 <= stage2_b_is_nan_10;
          stage2_exponent_09 <= stage2_exponent_10;
          stage2_zi_09 <= insn_o_1_819_0;
      end
      st_1_44 <= st_1_43;
      if (st_1_44) begin
          stage2_di_08 <= stage2_di_09;
          stage2_sign_08 <= stage2_sign_09;
          stage2_a_is_zero_08 <= stage2_a_is_zero_09;
          stage2_a_is_inf_08 <= stage2_a_is_inf_09;
          stage2_a_is_nan_08 <= stage2_a_is_nan_09;
          stage2_b_is_zero_08 <= stage2_b_is_zero_09;
          stage2_b_is_inf_08 <= stage2_b_is_inf_09;
          stage2_b_is_nan_08 <= stage2_b_is_nan_09;
          stage2_exponent_08 <= stage2_exponent_09;
          stage2_zi_08 <= insn_o_1_838_0;
      end
      st_1_45 <= st_1_44;
      if (st_1_45) begin
          stage2_di_07 <= stage2_di_08;
          stage2_sign_07 <= stage2_sign_08;
          stage2_a_is_zero_07 <= stage2_a_is_zero_08;
          stage2_a_is_inf_07 <= stage2_a_is_inf_08;
          stage2_a_is_nan_07 <= stage2_a_is_nan_08;
          stage2_b_is_zero_07 <= stage2_b_is_zero_08;
          stage2_b_is_inf_07 <= stage2_b_is_inf_08;
          stage2_b_is_nan_07 <= stage2_b_is_nan_08;
          stage2_exponent_07 <= stage2_exponent_08;
          stage2_zi_07 <= insn_o_1_857_0;
      end
      st_1_46 <= st_1_45;
      if (st_1_46) begin
          stage2_di_06 <= stage2_di_07;
          stage2_sign_06 <= stage2_sign_07;
          stage2_a_is_zero_06 <= stage2_a_is_zero_07;
          stage2_a_is_inf_06 <= stage2_a_is_inf_07;
          stage2_a_is_nan_06 <= stage2_a_is_nan_07;
          stage2_b_is_zero_06 <= stage2_b_is_zero_07;
          stage2_b_is_inf_06 <= stage2_b_is_inf_07;
          stage2_b_is_nan_06 <= stage2_b_is_nan_07;
          stage2_exponent_06 <= stage2_exponent_07;
          stage2_zi_06 <= insn_o_1_876_0;
      end
      st_1_47 <= st_1_46;
      if (st_1_47) begin
          stage2_di_05 <= stage2_di_06;
          stage2_sign_05 <= stage2_sign_06;
          stage2_a_is_zero_05 <= stage2_a_is_zero_06;
          stage2_a_is_inf_05 <= stage2_a_is_inf_06;
          stage2_a_is_nan_05 <= stage2_a_is_nan_06;
          stage2_b_is_zero_05 <= stage2_b_is_zero_06;
          stage2_b_is_inf_05 <= stage2_b_is_inf_06;
          stage2_b_is_nan_05 <= stage2_b_is_nan_06;
          stage2_exponent_05 <= stage2_exponent_06;
          stage2_zi_05 <= insn_o_1_895_0;
      end
      st_1_48 <= st_1_47;
      if (st_1_48) begin
          stage2_di_04 <= stage2_di_05;
          stage2_sign_04 <= stage2_sign_05;
          stage2_a_is_zero_04 <= stage2_a_is_zero_05;
          stage2_a_is_inf_04 <= stage2_a_is_inf_05;
          stage2_a_is_nan_04 <= stage2_a_is_nan_05;
          stage2_b_is_zero_04 <= stage2_b_is_zero_05;
          stage2_b_is_inf_04 <= stage2_b_is_inf_05;
          stage2_b_is_nan_04 <= stage2_b_is_nan_05;
          stage2_exponent_04 <= stage2_exponent_05;
          stage2_zi_04 <= insn_o_1_914_0;
      end
      st_1_49 <= st_1_48;
      if (st_1_49) begin
          stage2_di_03 <= stage2_di_04;
          stage2_sign_03 <= stage2_sign_04;
          stage2_a_is_zero_03 <= stage2_a_is_zero_04;
          stage2_a_is_inf_03 <= stage2_a_is_inf_04;
          stage2_a_is_nan_03 <= stage2_a_is_nan_04;
          stage2_b_is_zero_03 <= stage2_b_is_zero_04;
          stage2_b_is_inf_03 <= stage2_b_is_inf_04;
          stage2_b_is_nan_03 <= stage2_b_is_nan_04;
          stage2_exponent_03 <= stage2_exponent_04;
          stage2_zi_03 <= insn_o_1_933_0;
      end
      st_1_50 <= st_1_49;
      if (st_1_50) begin
          stage2_di_02 <= stage2_di_03;
          stage2_sign_02 <= stage2_sign_03;
          stage2_a_is_zero_02 <= stage2_a_is_zero_03;
          stage2_a_is_inf_02 <= stage2_a_is_inf_03;
          stage2_a_is_nan_02 <= stage2_a_is_nan_03;
          stage2_b_is_zero_02 <= stage2_b_is_zero_03;
          stage2_b_is_inf_02 <= stage2_b_is_inf_03;
          stage2_b_is_nan_02 <= stage2_b_is_nan_03;
          stage2_exponent_02 <= stage2_exponent_03;
          stage2_zi_02 <= insn_o_1_952_0;
      end
      st_1_51 <= st_1_50;
      if (st_1_51) begin
          stage2_di_01 <= stage2_di_02;
          stage2_sign_01 <= stage2_sign_02;
          stage2_a_is_zero_01 <= stage2_a_is_zero_02;
          stage2_a_is_inf_01 <= stage2_a_is_inf_02;
          stage2_a_is_nan_01 <= stage2_a_is_nan_02;
          stage2_b_is_zero_01 <= stage2_b_is_zero_02;
          stage2_b_is_inf_01 <= stage2_b_is_inf_02;
          stage2_b_is_nan_01 <= stage2_b_is_nan_02;
          stage2_exponent_01 <= stage2_exponent_02;
          stage2_zi_01 <= insn_o_1_971_0;
      end
      st_1_52 <= st_1_51;
      if (st_1_52) begin
          stage2_di_00 <= stage2_di_01;
          stage2_sign_00 <= stage2_sign_01;
          stage2_a_is_zero_00 <= stage2_a_is_zero_01;
          stage2_a_is_inf_00 <= stage2_a_is_inf_01;
          stage2_a_is_nan_00 <= stage2_a_is_nan_01;
          stage2_b_is_zero_00 <= stage2_b_is_zero_01;
          stage2_b_is_inf_00 <= stage2_b_is_inf_01;
          stage2_b_is_nan_00 <= stage2_b_is_nan_01;
          stage2_zi_00 <= insn_o_1_990_0;
          stage2_exponent_00 <= insn_o_1_999_0;
      end
      st_1_53 <= st_1_52;
      if (st_1_53) begin
          stage3_sign <= stage2_sign_00;
          stage3_a_is_zero <= stage2_a_is_zero_00;
          stage3_a_is_inf <= stage2_a_is_inf_00;
          stage3_a_is_nan <= stage2_a_is_nan_00;
          stage3_b_is_zero <= stage2_b_is_zero_00;
          stage3_b_is_inf <= stage2_b_is_inf_00;
          stage3_b_is_nan <= stage2_b_is_nan_00;
          stage3_fraction <= insn_o_1_1006_0;
          stage3_exponent <= insn_o_1_1008_0;
      end
      st_1_54 <= st_1_53;
      if (st_1_54) begin
          stage4_sign <= stage3_sign;
          stage4_a_is_zero <= stage3_a_is_zero;
          stage4_a_is_inf <= stage3_a_is_inf;
          stage4_a_is_nan <= stage3_a_is_nan;
          stage4_b_is_zero <= stage3_b_is_zero;
          stage4_b_is_inf <= stage3_b_is_inf;
          stage4_b_is_nan <= stage3_b_is_nan;
          stage4_fraction <= insn_o_1_1024_0;
          stage4_exponent <= insn_o_1_1027_0;
      end
      st_1_55 <= st_1_54;
      if (st_1_55) begin
          z_out <= stage5_result;
      end
    end
  end

endmodule
