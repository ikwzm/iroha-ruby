// Generated from iroha-0.1.0.

module fmul(clk, rst_n, i_valid, z_out, a_in, b_in);
  input clk;
  input rst_n;
  input i_valid;
  output [31:0] z_out;
  input [31:0] a_in;
  input [31:0] b_in;
  reg [31:0] z_out;

  // State decls
  reg st_1_1;
  reg st_1_2;
  reg st_1_3;
  reg st_1_4;
  reg st_1_5;
  // State vars
  // Registers
  wire  [0:0] start;
  reg  [23:0] stage1_a_fraction;
  reg  [7:0] stage1_a_exponent;
  reg  stage1_a_sign;
  reg  stage1_a_exponent_is_all_0;
  reg  stage1_a_fraction_is_all_0;
  reg  [23:0] stage1_b_fraction;
  reg  [7:0] stage1_b_exponent;
  reg  stage1_b_sign;
  reg  stage1_b_exponent_is_all_0;
  reg  stage1_b_fraction_is_all_0;
  reg  [47:0] stage2_fraction;
  reg  signed [9:0] stage2_exponent;
  reg  stage2_sign;
  reg  stage2_a_is_zero;
  reg  stage2_a_is_inf;
  reg  stage2_a_is_nan;
  reg  stage2_b_is_zero;
  reg  stage2_b_is_inf;
  reg  stage2_b_is_nan;
  reg  [22:0] stage3_fraction;
  reg  signed [9:0] stage3_exponent;
  reg  stage3_sign;
  reg  stage3_guard;
  reg  stage3_round;
  reg  stage3_sticky;
  reg  stage3_a_is_zero;
  reg  stage3_a_is_inf;
  reg  stage3_a_is_nan;
  reg  stage3_b_is_zero;
  reg  stage3_b_is_inf;
  reg  stage3_b_is_nan;
  reg  [22:0] stage4_fraction;
  reg  signed [9:0] stage4_exponent;
  reg  stage4_sign;
  reg  stage4_a_is_zero;
  reg  stage4_a_is_inf;
  reg  stage4_a_is_nan;
  reg  stage4_b_is_zero;
  reg  stage4_b_is_inf;
  reg  stage4_b_is_nan;
  wire  [31:0] stage1_a_data_in;
  wire  [7:0] stage1_a_exponent_in;
  wire  [22:0] stage1_a_fraction_in;
  wire  stage1_a_sign_in;
  wire  stage1_a_exponent_zero;
  wire  [0:0] stage1_a_fraction_msb;
  wire  [31:0] stage1_b_data_in;
  wire  [7:0] stage1_b_exponent_in;
  wire  [22:0] stage1_b_fraction_in;
  wire  stage1_b_sign_in;
  wire  stage1_b_exponent_zero;
  wire  [0:0] stage1_b_fraction_msb;
  wire  [9:0] stage2_exponent_a_in;
  wire  signed [9:0] stage2_exponent_a_d;
  wire  [9:0] stage2_exponent_b_in;
  wire  signed [9:0] stage2_exponent_b_d;
  wire  stage2_exponent_a_is_all_0;
  wire  stage2_exponent_a_is_all_1;
  wire  stage2_fraction_a_is_all_0;
  wire  stage2_fraction_a_is_not_0;
  wire  stage2_exponent_b_is_all_0;
  wire  stage2_exponent_b_is_all_1;
  wire  stage2_fraction_b_is_all_0;
  wire  stage2_fraction_b_is_not_0;
  wire  [0:0] stage3_mul_fraction_msb;
  wire  signed [9:0] stage3_mul_exponent;
  wire  [22:0] stage3_mul_0_fraction;
  wire  stage3_mul_0_guard;
  wire  stage3_mul_0_round;
  wire  stage3_mul_0_sticky;
  wire  [20:0] stage3_mul_0_sticky_data;
  wire  anon_103;
  wire  [22:0] stage3_mul_1_fraction;
  wire  stage3_mul_1_guard;
  wire  stage3_mul_1_round;
  wire  stage3_mul_1_sticky;
  wire  [21:0] stage3_mul_1_sticky_data;
  wire  anon_116;
  wire  stage4_fraction_lsb;
  wire  [0:0] stage4_fraction_increment;
  wire  anon_120;
  wire  anon_121;
  wire  [0:0] stage4_exponent_increment;
  wire  anon_124;
  wire  stage5_exp_natural;
  wire  stage5_exp_underflow;
  wire  stage5_exp_overflow;
  wire  [7:0] stage5_exponent_in;
  wire  [22:0] stage5_fraction_in;
  wire  [7:0] stage5_exponent_i1;
  wire  [22:0] stage5_fraction_i1;
  wire  [7:0] stage5_exponent_di;
  wire  [22:0] stage5_fraction_di;
  wire  stage5_a_is_zero;
  wire  stage5_a_is_inf;
  wire  stage5_a_is_nan;
  wire  stage5_a_is_norm;
  wire  anon_150;
  wire  anon_151;
  wire  stage5_b_is_zero;
  wire  stage5_b_is_inf;
  wire  stage5_b_is_nan;
  wire  stage5_b_is_norm;
  wire  anon_156;
  wire  anon_157;
  wire  stage5_set_zero;
  wire  anon_159;
  wire  anon_160;
  wire  anon_161;
  wire  anon_162;
  wire  stage5_set_inf;
  wire  anon_164;
  wire  anon_165;
  wire  anon_166;
  wire  anon_167;
  wire  stage5_set_norm;
  wire  stage5_set_nan;
  wire  [22:0] stage5_fraction_o0;
  wire  [7:0] stage5_exponent_o0;
  wire  [22:0] stage5_fraction_o1;
  wire  [7:0] stage5_exponent_o1;
  wire  [0:0] stage5_sign_o;
  wire  [22:0] stage5_fraction_o;
  wire  [7:0] stage5_exponent_o;
  wire  [31:0] stage5_result;
  // Resources
  // eq:10
  wire [7:0] eq_10_s0;
  assign eq_10_s0 = stage1_a_exponent_in;
  wire [7:0] eq_10_s1;
  assign eq_10_s1 = 8'd0;
  wire eq_10_d0;
  assign eq_10_d0 = eq_10_s0 == eq_10_s1;
  // eq:16
  wire [22:0] eq_16_s0;
  assign eq_16_s0 = stage1_a_fraction_in;
  wire [22:0] eq_16_s1;
  assign eq_16_s1 = 23'd0;
  wire eq_16_d0;
  assign eq_16_d0 = eq_16_s0 == eq_16_s1;
  // eq:20
  wire [7:0] eq_20_s0;
  assign eq_20_s0 = stage1_b_exponent_in;
  wire [7:0] eq_20_s1;
  assign eq_20_s1 = 8'd0;
  wire eq_20_d0;
  assign eq_20_d0 = eq_20_s0 == eq_20_s1;
  // eq:26
  wire [22:0] eq_26_s0;
  assign eq_26_s0 = stage1_b_fraction_in;
  wire [22:0] eq_26_s1;
  assign eq_26_s1 = 23'd0;
  wire eq_26_d0;
  assign eq_26_d0 = eq_26_s0 == eq_26_s1;
  // sub:28
  wire [9:0] sub_28_s0;
  assign sub_28_s0 = stage2_exponent_a_in;
  wire [7:0] sub_28_s1;
  assign sub_28_s1 = 8'd127;
  wire signed [9:0] sub_28_d0;
  assign sub_28_d0 = sub_28_s0 - sub_28_s1;
  // sub:30
  wire [9:0] sub_30_s0;
  assign sub_30_s0 = stage2_exponent_b_in;
  wire [7:0] sub_30_s1;
  assign sub_30_s1 = 8'd127;
  wire signed [9:0] sub_30_d0;
  assign sub_30_d0 = sub_30_s0 - sub_30_s1;
  // add:31
  wire signed [9:0] add_31_s0;
  assign add_31_s0 = stage2_exponent_a_d;
  wire signed [9:0] add_31_s1;
  assign add_31_s1 = stage2_exponent_b_d;
  wire signed [9:0] add_31_d0;
  assign add_31_d0 = add_31_s0 + add_31_s1;
  // mul:32
  wire [23:0] mul_32_s0;
  assign mul_32_s0 = stage1_a_fraction;
  wire [23:0] mul_32_s1;
  assign mul_32_s1 = stage1_b_fraction;
  wire [47:0] mul_32_d0;
  assign mul_32_d0 = mul_32_s0 * mul_32_s1;
  // eq:35
  wire [7:0] eq_35_s0;
  assign eq_35_s0 = stage1_a_exponent;
  wire [7:0] eq_35_s1;
  assign eq_35_s1 = 8'd255;
  wire eq_35_d0;
  assign eq_35_d0 = eq_35_s0 == eq_35_s1;
  // eq:42
  wire [7:0] eq_42_s0;
  assign eq_42_s0 = stage1_b_exponent;
  wire [7:0] eq_42_s1;
  assign eq_42_s1 = 8'd255;
  wire eq_42_d0;
  assign eq_42_d0 = eq_42_s0 == eq_42_s1;
  // add:49
  wire signed [9:0] add_49_s0;
  assign add_49_s0 = stage2_exponent;
  wire [0:0] add_49_s1;
  assign add_49_s1 = stage3_mul_fraction_msb;
  wire signed [9:0] add_49_d0;
  assign add_49_d0 = add_49_s0 + add_49_s1;
  // eq:54
  wire [20:0] eq_54_s0;
  assign eq_54_s0 = stage3_mul_0_sticky_data;
  wire [20:0] eq_54_s1;
  assign eq_54_s1 = 21'd0;
  wire eq_54_d0;
  assign eq_54_d0 = eq_54_s0 == eq_54_s1;
  // eq:60
  wire [21:0] eq_60_s0;
  assign eq_60_s0 = stage3_mul_1_sticky_data;
  wire [21:0] eq_60_s1;
  assign eq_60_s1 = 22'd0;
  wire eq_60_d0;
  assign eq_60_d0 = eq_60_s0 == eq_60_s1;
  // add:62
  wire signed [9:0] add_62_s0;
  assign add_62_s0 = stage3_mul_exponent;
  wire [7:0] add_62_s1;
  assign add_62_s1 = 8'd127;
  wire signed [9:0] add_62_d0;
  assign add_62_d0 = add_62_s0 + add_62_s1;
  // eq:78
  wire [22:0] eq_78_s0;
  assign eq_78_s0 = stage3_fraction;
  wire [22:0] eq_78_s1;
  assign eq_78_s1 = 23'd8388607;
  wire eq_78_d0;
  assign eq_78_d0 = eq_78_s0 == eq_78_s1;
  // add:80
  wire [22:0] add_80_s0;
  assign add_80_s0 = stage3_fraction;
  wire [0:0] add_80_s1;
  assign add_80_s1 = stage4_fraction_increment;
  wire [22:0] add_80_d0;
  assign add_80_d0 = add_80_s0 + add_80_s1;
  // add:81
  wire signed [9:0] add_81_s0;
  assign add_81_s0 = stage3_exponent;
  wire [0:0] add_81_s1;
  assign add_81_s1 = stage4_exponent_increment;
  wire signed [9:0] add_81_d0;
  assign add_81_d0 = add_81_s0 + add_81_s1;
  // gt:89
  wire signed [9:0] gt_89_s0;
  assign gt_89_s0 = stage4_exponent;
  wire signed [9:0] gt_89_s1;
  assign gt_89_s1 = 10'd0;
  wire gt_89_d0;
  assign gt_89_d0 = gt_89_s0 > gt_89_s1;
  // gte:91
  wire signed [9:0] gte_91_s0;
  assign gte_91_s0 = stage4_exponent;
  wire signed [9:0] gte_91_s1;
  assign gte_91_s1 = 10'd255;
  wire gte_91_d0;
  assign gte_91_d0 = gte_91_s0 >= gte_91_s1;
  // Insn wires
  wire  [0:0] insn_o_1_6_0;
  wire  [31:0] insn_o_1_7_0;
  wire  [7:0] insn_o_1_8_0;
  wire  [22:0] insn_o_1_9_0;
  wire  insn_o_1_10_0;
  wire  insn_o_1_11_0;
  wire  [0:0] insn_o_1_12_0;
  wire  [23:0] insn_o_1_13_0;
  wire  [7:0] insn_o_1_14_0;
  wire  insn_o_1_15_0;
  wire  insn_o_1_16_0;
  wire  insn_o_1_17_0;
  wire  [31:0] insn_o_1_18_0;
  wire  [7:0] insn_o_1_19_0;
  wire  [22:0] insn_o_1_20_0;
  wire  insn_o_1_21_0;
  wire  insn_o_1_22_0;
  wire  [0:0] insn_o_1_23_0;
  wire  [23:0] insn_o_1_24_0;
  wire  [7:0] insn_o_1_25_0;
  wire  insn_o_1_26_0;
  wire  insn_o_1_27_0;
  wire  insn_o_1_28_0;
  wire  [9:0] insn_o_1_30_0;
  wire  signed [9:0] insn_o_1_31_0;
  wire  [9:0] insn_o_1_32_0;
  wire  signed [9:0] insn_o_1_33_0;
  wire  signed [9:0] insn_o_1_34_0;
  wire  [47:0] insn_o_1_35_0;
  wire  insn_o_1_36_0;
  wire  insn_o_1_37_0;
  wire  insn_o_1_38_0;
  wire  insn_o_1_39_0;
  wire  insn_o_1_40_0;
  wire  insn_o_1_41_0;
  wire  insn_o_1_42_0;
  wire  insn_o_1_43_0;
  wire  insn_o_1_44_0;
  wire  insn_o_1_45_0;
  wire  insn_o_1_46_0;
  wire  insn_o_1_47_0;
  wire  insn_o_1_48_0;
  wire  insn_o_1_49_0;
  wire  insn_o_1_50_0;
  wire  [0:0] insn_o_1_52_0;
  wire  signed [9:0] insn_o_1_53_0;
  wire  [22:0] insn_o_1_54_0;
  wire  insn_o_1_55_0;
  wire  insn_o_1_56_0;
  wire  [20:0] insn_o_1_57_0;
  wire  insn_o_1_58_0;
  wire  insn_o_1_59_0;
  wire  [22:0] insn_o_1_60_0;
  wire  insn_o_1_61_0;
  wire  insn_o_1_62_0;
  wire  [21:0] insn_o_1_63_0;
  wire  insn_o_1_64_0;
  wire  insn_o_1_65_0;
  wire  signed [9:0] insn_o_1_66_0;
  wire  [22:0] insn_o_1_67_0;
  wire  insn_o_1_68_0;
  wire  insn_o_1_69_0;
  wire  insn_o_1_70_0;
  wire  insn_o_1_71_0;
  wire  insn_o_1_72_0;
  wire  insn_o_1_73_0;
  wire  insn_o_1_74_0;
  wire  insn_o_1_75_0;
  wire  insn_o_1_76_0;
  wire  insn_o_1_77_0;
  wire  insn_o_1_79_0;
  wire  insn_o_1_80_0;
  wire  insn_o_1_81_0;
  wire  [0:0] insn_o_1_82_0;
  wire  insn_o_1_83_0;
  wire  [0:0] insn_o_1_84_0;
  wire  [22:0] insn_o_1_85_0;
  wire  signed [9:0] insn_o_1_86_0;
  wire  insn_o_1_87_0;
  wire  insn_o_1_88_0;
  wire  insn_o_1_89_0;
  wire  insn_o_1_90_0;
  wire  insn_o_1_91_0;
  wire  insn_o_1_92_0;
  wire  insn_o_1_93_0;
  wire  insn_o_1_95_0;
  wire  insn_o_1_96_0;
  wire  insn_o_1_97_0;
  wire  [7:0] insn_o_1_98_0;
  wire  [22:0] insn_o_1_99_0;
  wire  [7:0] insn_o_1_100_0;
  wire  [22:0] insn_o_1_101_0;
  wire  [7:0] insn_o_1_102_0;
  wire  [22:0] insn_o_1_103_0;
  wire  insn_o_1_104_0;
  wire  insn_o_1_105_0;
  wire  insn_o_1_106_0;
  wire  insn_o_1_107_0;
  wire  insn_o_1_108_0;
  wire  insn_o_1_109_0;
  wire  insn_o_1_110_0;
  wire  insn_o_1_111_0;
  wire  insn_o_1_112_0;
  wire  insn_o_1_113_0;
  wire  insn_o_1_114_0;
  wire  insn_o_1_115_0;
  wire  insn_o_1_116_0;
  wire  insn_o_1_117_0;
  wire  insn_o_1_118_0;
  wire  insn_o_1_119_0;
  wire  insn_o_1_120_0;
  wire  insn_o_1_121_0;
  wire  insn_o_1_122_0;
  wire  insn_o_1_123_0;
  wire  insn_o_1_124_0;
  wire  insn_o_1_125_0;
  wire  insn_o_1_126_0;
  wire  insn_o_1_127_0;
  wire  [22:0] insn_o_1_128_0;
  wire  [7:0] insn_o_1_129_0;
  wire  [22:0] insn_o_1_130_0;
  wire  [7:0] insn_o_1_131_0;
  wire  [0:0] insn_o_1_132_0;
  wire  [22:0] insn_o_1_133_0;
  wire  [7:0] insn_o_1_134_0;
  wire  [31:0] insn_o_1_135_0;
  // Insn assigns
  assign insn_o_1_6_0 = i_valid;
  assign start = insn_o_1_6_0;
  assign insn_o_1_7_0 = a_in;
  assign stage1_a_data_in = insn_o_1_7_0;
  assign insn_o_1_8_0 = stage1_a_data_in[30:23];
  assign stage1_a_exponent_in = insn_o_1_8_0;
  assign insn_o_1_9_0 = stage1_a_data_in[22:0];
  assign stage1_a_fraction_in = insn_o_1_9_0;
  assign insn_o_1_10_0 = stage1_a_data_in[31:31];
  assign stage1_a_sign_in = insn_o_1_10_0;
  assign insn_o_1_11_0 = eq_10_d0;
  assign stage1_a_exponent_zero = insn_o_1_11_0;
  assign insn_o_1_12_0 = ~stage1_a_exponent_zero;
  assign stage1_a_fraction_msb = insn_o_1_12_0;
  assign insn_o_1_13_0 = {stage1_a_fraction_msb, stage1_a_fraction_in};
  assign insn_o_1_17_0 = eq_16_d0;
  assign insn_o_1_18_0 = b_in;
  assign stage1_b_data_in = insn_o_1_18_0;
  assign insn_o_1_19_0 = stage1_b_data_in[30:23];
  assign stage1_b_exponent_in = insn_o_1_19_0;
  assign insn_o_1_20_0 = stage1_b_data_in[22:0];
  assign stage1_b_fraction_in = insn_o_1_20_0;
  assign insn_o_1_21_0 = stage1_b_data_in[31:31];
  assign stage1_b_sign_in = insn_o_1_21_0;
  assign insn_o_1_22_0 = eq_20_d0;
  assign stage1_b_exponent_zero = insn_o_1_22_0;
  assign insn_o_1_23_0 = ~stage1_b_exponent_zero;
  assign stage1_b_fraction_msb = insn_o_1_23_0;
  assign insn_o_1_24_0 = {stage1_b_fraction_msb, stage1_b_fraction_in};
  assign insn_o_1_28_0 = eq_26_d0;
  assign insn_o_1_30_0 = {2'd0, stage1_a_exponent};
  assign stage2_exponent_a_in = insn_o_1_30_0;
  assign insn_o_1_31_0 = sub_28_d0;
  assign stage2_exponent_a_d = insn_o_1_31_0;
  assign insn_o_1_32_0 = {2'd0, stage1_b_exponent};
  assign stage2_exponent_b_in = insn_o_1_32_0;
  assign insn_o_1_33_0 = sub_30_d0;
  assign stage2_exponent_b_d = insn_o_1_33_0;
  assign insn_o_1_34_0 = add_31_d0;
  assign insn_o_1_35_0 = mul_32_d0;
  assign insn_o_1_36_0 = stage1_a_sign ^ stage1_b_sign;
  assign stage2_exponent_a_is_all_0 = stage1_a_exponent_is_all_0;
  assign insn_o_1_38_0 = eq_35_d0;
  assign stage2_exponent_a_is_all_1 = insn_o_1_38_0;
  assign stage2_fraction_a_is_all_0 = stage1_a_fraction_is_all_0;
  assign insn_o_1_40_0 = ~stage1_a_fraction_is_all_0;
  assign stage2_fraction_a_is_not_0 = insn_o_1_40_0;
  assign insn_o_1_41_0 = stage2_exponent_a_is_all_0 & stage2_fraction_a_is_all_0;
  assign insn_o_1_42_0 = stage2_exponent_a_is_all_1 & stage2_fraction_a_is_all_0;
  assign insn_o_1_43_0 = stage2_exponent_a_is_all_1 & stage2_fraction_a_is_not_0;
  assign stage2_exponent_b_is_all_0 = stage1_b_exponent_is_all_0;
  assign insn_o_1_45_0 = eq_42_d0;
  assign stage2_exponent_b_is_all_1 = insn_o_1_45_0;
  assign stage2_fraction_b_is_all_0 = stage1_b_fraction_is_all_0;
  assign insn_o_1_47_0 = ~stage1_b_fraction_is_all_0;
  assign stage2_fraction_b_is_not_0 = insn_o_1_47_0;
  assign insn_o_1_48_0 = stage2_exponent_b_is_all_0 & stage2_fraction_b_is_all_0;
  assign insn_o_1_49_0 = stage2_exponent_b_is_all_1 & stage2_fraction_b_is_all_0;
  assign insn_o_1_50_0 = stage2_exponent_b_is_all_1 & stage2_fraction_b_is_not_0;
  assign insn_o_1_52_0 = stage2_fraction[47:47];
  assign stage3_mul_fraction_msb = insn_o_1_52_0;
  assign insn_o_1_53_0 = add_49_d0;
  assign stage3_mul_exponent = insn_o_1_53_0;
  assign insn_o_1_54_0 = stage2_fraction[45:23];
  assign stage3_mul_0_fraction = insn_o_1_54_0;
  assign insn_o_1_55_0 = stage2_fraction[22:22];
  assign stage3_mul_0_guard = insn_o_1_55_0;
  assign insn_o_1_56_0 = stage2_fraction[21:21];
  assign stage3_mul_0_round = insn_o_1_56_0;
  assign insn_o_1_57_0 = stage2_fraction[20:0];
  assign stage3_mul_0_sticky_data = insn_o_1_57_0;
  assign insn_o_1_58_0 = eq_54_d0;
  assign anon_103 = insn_o_1_58_0;
  assign insn_o_1_59_0 = ~anon_103;
  assign stage3_mul_0_sticky = insn_o_1_59_0;
  assign insn_o_1_60_0 = stage2_fraction[46:24];
  assign stage3_mul_1_fraction = insn_o_1_60_0;
  assign insn_o_1_61_0 = stage2_fraction[23:23];
  assign stage3_mul_1_guard = insn_o_1_61_0;
  assign insn_o_1_62_0 = stage2_fraction[22:22];
  assign stage3_mul_1_round = insn_o_1_62_0;
  assign insn_o_1_63_0 = stage2_fraction[21:0];
  assign stage3_mul_1_sticky_data = insn_o_1_63_0;
  assign insn_o_1_64_0 = eq_60_d0;
  assign anon_116 = insn_o_1_64_0;
  assign insn_o_1_65_0 = ~anon_116;
  assign stage3_mul_1_sticky = insn_o_1_65_0;
  assign insn_o_1_66_0 = add_62_d0;
  assign insn_o_1_67_0 = stage3_mul_fraction_msb ? stage3_mul_1_fraction : stage3_mul_0_fraction;
  assign insn_o_1_68_0 = stage3_mul_fraction_msb ? stage3_mul_1_guard : stage3_mul_0_guard;
  assign insn_o_1_69_0 = stage3_mul_fraction_msb ? stage3_mul_1_round : stage3_mul_0_round;
  assign insn_o_1_70_0 = stage3_mul_fraction_msb ? stage3_mul_1_sticky : stage3_mul_0_sticky;
  assign insn_o_1_79_0 = stage3_fraction[0:0];
  assign stage4_fraction_lsb = insn_o_1_79_0;
  assign insn_o_1_80_0 = stage4_fraction_lsb | stage3_round;
  assign anon_120 = insn_o_1_80_0;
  assign insn_o_1_81_0 = anon_120 | stage3_sticky;
  assign anon_121 = insn_o_1_81_0;
  assign insn_o_1_82_0 = stage3_guard & anon_121;
  assign stage4_fraction_increment = insn_o_1_82_0;
  assign insn_o_1_83_0 = eq_78_d0;
  assign anon_124 = insn_o_1_83_0;
  assign insn_o_1_84_0 = stage4_fraction_increment & anon_124;
  assign stage4_exponent_increment = insn_o_1_84_0;
  assign insn_o_1_85_0 = add_80_d0;
  assign insn_o_1_86_0 = add_81_d0;
  assign insn_o_1_95_0 = gt_89_d0;
  assign stage5_exp_natural = insn_o_1_95_0;
  assign insn_o_1_96_0 = ~stage5_exp_natural;
  assign stage5_exp_underflow = insn_o_1_96_0;
  assign insn_o_1_97_0 = gte_91_d0;
  assign stage5_exp_overflow = insn_o_1_97_0;
  assign insn_o_1_98_0 = stage4_exponent[7:0];
  assign stage5_exponent_in = insn_o_1_98_0;
  assign stage5_fraction_in = stage4_fraction;
  assign insn_o_1_100_0 = stage5_exp_overflow ? 8'd255 : stage5_exponent_in;
  assign stage5_exponent_i1 = insn_o_1_100_0;
  assign insn_o_1_101_0 = stage5_exp_overflow ? 23'd0 : stage5_fraction_in;
  assign stage5_fraction_i1 = insn_o_1_101_0;
  assign insn_o_1_102_0 = stage5_exp_underflow ? 8'd0 : stage5_exponent_i1;
  assign stage5_exponent_di = insn_o_1_102_0;
  assign insn_o_1_103_0 = stage5_exp_underflow ? 23'd0 : stage5_fraction_i1;
  assign stage5_fraction_di = insn_o_1_103_0;
  assign stage5_a_is_zero = stage4_a_is_zero;
  assign stage5_a_is_inf = stage4_a_is_inf;
  assign stage5_a_is_nan = stage4_a_is_nan;
  assign insn_o_1_107_0 = stage5_a_is_zero | stage5_a_is_inf;
  assign anon_150 = insn_o_1_107_0;
  assign insn_o_1_108_0 = anon_150 | stage5_a_is_nan;
  assign anon_151 = insn_o_1_108_0;
  assign insn_o_1_109_0 = ~anon_151;
  assign stage5_a_is_norm = insn_o_1_109_0;
  assign stage5_b_is_zero = stage4_b_is_zero;
  assign stage5_b_is_inf = stage4_b_is_inf;
  assign stage5_b_is_nan = stage4_b_is_nan;
  assign insn_o_1_113_0 = stage5_b_is_zero | stage5_b_is_inf;
  assign anon_156 = insn_o_1_113_0;
  assign insn_o_1_114_0 = anon_156 | stage5_b_is_nan;
  assign anon_157 = insn_o_1_114_0;
  assign insn_o_1_115_0 = ~anon_157;
  assign stage5_b_is_norm = insn_o_1_115_0;
  assign insn_o_1_116_0 = stage5_a_is_zero & stage5_b_is_zero;
  assign anon_159 = insn_o_1_116_0;
  assign insn_o_1_117_0 = stage5_a_is_zero & stage5_b_is_norm;
  assign anon_160 = insn_o_1_117_0;
  assign insn_o_1_118_0 = anon_159 | anon_160;
  assign anon_161 = insn_o_1_118_0;
  assign insn_o_1_119_0 = stage5_a_is_norm & stage5_b_is_zero;
  assign anon_162 = insn_o_1_119_0;
  assign insn_o_1_120_0 = anon_161 | anon_162;
  assign stage5_set_zero = insn_o_1_120_0;
  assign insn_o_1_121_0 = stage5_a_is_inf & stage5_b_is_inf;
  assign anon_164 = insn_o_1_121_0;
  assign insn_o_1_122_0 = stage5_a_is_inf & stage5_b_is_norm;
  assign anon_165 = insn_o_1_122_0;
  assign insn_o_1_123_0 = anon_164 | anon_165;
  assign anon_166 = insn_o_1_123_0;
  assign insn_o_1_124_0 = stage5_a_is_norm & stage5_b_is_inf;
  assign anon_167 = insn_o_1_124_0;
  assign insn_o_1_125_0 = anon_166 | anon_167;
  assign stage5_set_inf = insn_o_1_125_0;
  assign insn_o_1_126_0 = stage5_a_is_norm & stage5_b_is_norm;
  assign stage5_set_norm = insn_o_1_126_0;
  assign insn_o_1_127_0 = stage5_a_is_nan | stage5_b_is_nan;
  assign stage5_set_nan = insn_o_1_127_0;
  assign insn_o_1_128_0 = stage5_set_norm ? stage5_fraction_di : 23'd2097152;
  assign stage5_fraction_o0 = insn_o_1_128_0;
  assign insn_o_1_129_0 = stage5_set_norm ? stage5_exponent_di : 8'd255;
  assign stage5_exponent_o0 = insn_o_1_129_0;
  assign insn_o_1_130_0 = stage5_set_inf ? 23'd0 : stage5_fraction_o0;
  assign stage5_fraction_o1 = insn_o_1_130_0;
  assign insn_o_1_131_0 = stage5_set_inf ? 8'd255 : stage5_exponent_o0;
  assign stage5_exponent_o1 = insn_o_1_131_0;
  assign insn_o_1_132_0 = stage5_set_nan ? 1'd0 : stage4_sign;
  assign stage5_sign_o = insn_o_1_132_0;
  assign insn_o_1_133_0 = stage5_set_zero ? 23'd0 : stage5_fraction_o1;
  assign stage5_fraction_o = insn_o_1_133_0;
  assign insn_o_1_134_0 = stage5_set_zero ? 8'd0 : stage5_exponent_o1;
  assign stage5_exponent_o = insn_o_1_134_0;
  assign insn_o_1_135_0 = {stage5_sign_o, stage5_exponent_o, stage5_fraction_o};
  assign stage5_result = insn_o_1_135_0;

  // Table 1
  always @(posedge clk) begin
    if (!rst_n) begin
      st_1_1 <= 0;
      st_1_2 <= 0;
      st_1_3 <= 0;
      st_1_4 <= 0;
      st_1_5 <= 0;
    end else begin
      if (start) begin
          stage1_a_exponent <= stage1_a_exponent_in;
          stage1_a_sign <= stage1_a_sign_in;
          stage1_a_exponent_is_all_0 <= stage1_a_exponent_zero;
          stage1_b_exponent <= stage1_b_exponent_in;
          stage1_b_sign <= stage1_b_sign_in;
          stage1_b_exponent_is_all_0 <= stage1_b_exponent_zero;
          stage1_a_fraction <= insn_o_1_13_0;
          stage1_a_fraction_is_all_0 <= insn_o_1_17_0;
          stage1_b_fraction <= insn_o_1_24_0;
          stage1_b_fraction_is_all_0 <= insn_o_1_28_0;
      end
      st_1_2 <= start;
      if (st_1_2) begin
          stage2_exponent <= insn_o_1_34_0;
          stage2_fraction <= insn_o_1_35_0;
          stage2_sign <= insn_o_1_36_0;
          stage2_a_is_zero <= insn_o_1_41_0;
          stage2_a_is_inf <= insn_o_1_42_0;
          stage2_a_is_nan <= insn_o_1_43_0;
          stage2_b_is_zero <= insn_o_1_48_0;
          stage2_b_is_inf <= insn_o_1_49_0;
          stage2_b_is_nan <= insn_o_1_50_0;
      end
      st_1_3 <= st_1_2;
      if (st_1_3) begin
          stage3_sign <= stage2_sign;
          stage3_a_is_zero <= stage2_a_is_zero;
          stage3_a_is_inf <= stage2_a_is_inf;
          stage3_a_is_nan <= stage2_a_is_nan;
          stage3_b_is_zero <= stage2_b_is_zero;
          stage3_b_is_inf <= stage2_b_is_inf;
          stage3_b_is_nan <= stage2_b_is_nan;
          stage3_exponent <= insn_o_1_66_0;
          stage3_fraction <= insn_o_1_67_0;
          stage3_guard <= insn_o_1_68_0;
          stage3_round <= insn_o_1_69_0;
          stage3_sticky <= insn_o_1_70_0;
      end
      st_1_4 <= st_1_3;
      if (st_1_4) begin
          stage4_sign <= stage3_sign;
          stage4_a_is_zero <= stage3_a_is_zero;
          stage4_a_is_inf <= stage3_a_is_inf;
          stage4_a_is_nan <= stage3_a_is_nan;
          stage4_b_is_zero <= stage3_b_is_zero;
          stage4_b_is_inf <= stage3_b_is_inf;
          stage4_b_is_nan <= stage3_b_is_nan;
          stage4_fraction <= insn_o_1_85_0;
          stage4_exponent <= insn_o_1_86_0;
      end
      st_1_5 <= st_1_4;
      if (st_1_5) begin
          z_out <= stage5_result;
      end
    end
  end

endmodule
